module control  (
	input  clock, reset,
	input  logic [11:0] in,
	output logic [11:0] out [148:0]
);
	logic [11:0] registers [148:0];
	assign out[0] = registers[0];
	assign out[1] = registers[1];
	assign out[2] = registers[2];
	assign out[3] = registers[3];
	assign out[4] = registers[4];
	assign out[5] = registers[5];
	assign out[6] = registers[6];
	assign out[7] = registers[7];
	assign out[8] = registers[8];
	assign out[9] = registers[9];
	assign out[10] = registers[10];
	assign out[11] = registers[11];
	assign out[12] = registers[12];
	assign out[13] = registers[13];
	assign out[14] = registers[14];
	assign out[15] = registers[15];
	assign out[16] = registers[16];
	assign out[17] = registers[17];
	assign out[18] = registers[18];
	assign out[19] = registers[19];
	assign out[20] = registers[20];
	assign out[21] = registers[21];
	assign out[22] = registers[22];
	assign out[23] = registers[23];
	assign out[24] = registers[24];
	assign out[25] = registers[25];
	assign out[26] = registers[26];
	assign out[27] = registers[27];
	assign out[28] = registers[28];
	assign out[29] = registers[29];
	assign out[30] = registers[30];
	assign out[31] = registers[31];
	assign out[32] = registers[32];
	assign out[33] = registers[33];
	assign out[34] = registers[34];
	assign out[35] = registers[35];
	assign out[36] = registers[36];
	assign out[37] = registers[37];
	assign out[38] = registers[38];
	assign out[39] = registers[39];
	assign out[40] = registers[40];
	assign out[41] = registers[41];
	assign out[42] = registers[42];
	assign out[43] = registers[43];
	assign out[44] = registers[44];
	assign out[45] = registers[45];
	assign out[46] = registers[46];
	assign out[47] = registers[47];
	assign out[48] = registers[48];
	assign out[49] = registers[49];
	assign out[50] = registers[50];
	assign out[51] = registers[51];
	assign out[52] = registers[52];
	assign out[53] = registers[53];
	assign out[54] = registers[54];
	assign out[55] = registers[55];
	assign out[56] = registers[56];
	assign out[57] = registers[57];
	assign out[58] = registers[58];
	assign out[59] = registers[59];
	assign out[60] = registers[60];
	assign out[61] = registers[61];
	assign out[62] = registers[62];
	assign out[63] = registers[63];
	assign out[64] = registers[64];
	assign out[65] = registers[65];
	assign out[66] = registers[66];
	assign out[67] = registers[67];
	assign out[68] = registers[68];
	assign out[69] = registers[69];
	assign out[70] = registers[70];
	assign out[71] = registers[71];
	assign out[72] = registers[72];
	assign out[73] = registers[73];
	assign out[74] = registers[74];
	assign out[75] = registers[75];
	assign out[76] = registers[76];
	assign out[77] = registers[77];
	assign out[78] = registers[78];
	assign out[79] = registers[79];
	assign out[80] = registers[80];
	assign out[81] = registers[81];
	assign out[82] = registers[82];
	assign out[83] = registers[83];
	assign out[84] = registers[84];
	assign out[85] = registers[85];
	assign out[86] = registers[86];
	assign out[87] = registers[87];
	assign out[88] = registers[88];
	assign out[89] = registers[89];
	assign out[90] = registers[90];
	assign out[91] = registers[91];
	assign out[92] = registers[92];
	assign out[93] = registers[93];
	assign out[94] = registers[94];
	assign out[95] = registers[95];
	assign out[96] = registers[96];
	assign out[97] = registers[97];
	assign out[98] = registers[98];
	assign out[99] = registers[99];
	assign out[100] = registers[100];
	assign out[101] = registers[101];
	assign out[102] = registers[102];
	assign out[103] = registers[103];
	assign out[104] = registers[104];
	assign out[105] = registers[105];
	assign out[106] = registers[106];
	assign out[107] = registers[107];
	assign out[108] = registers[108];
	assign out[109] = registers[109];
	assign out[110] = registers[110];
	assign out[111] = registers[111];
	assign out[112] = registers[112];
	assign out[113] = registers[113];
	assign out[114] = registers[114];
	assign out[115] = registers[115];
	assign out[116] = registers[116];
	assign out[117] = registers[117];
	assign out[118] = registers[118];
	assign out[119] = registers[119];
	assign out[120] = registers[120];
	assign out[121] = registers[121];
	assign out[122] = registers[122];
	assign out[123] = registers[123];
	assign out[124] = registers[124];
	assign out[125] = registers[125];
	assign out[126] = registers[126];
	assign out[127] = registers[127];
	assign out[128] = registers[128];
	assign out[129] = registers[129];
	assign out[130] = registers[130];
	assign out[131] = registers[131];
	assign out[132] = registers[132];
	assign out[133] = registers[133];
	assign out[134] = registers[134];
	assign out[135] = registers[135];
	assign out[136] = registers[136];
	assign out[137] = registers[137];
	assign out[138] = registers[138];
	assign out[139] = registers[139];
	assign out[140] = registers[140];
	assign out[141] = registers[141];
	assign out[142] = registers[142];
	assign out[143] = registers[143];
	assign out[144] = registers[144];
	assign out[145] = registers[145];
	assign out[146] = registers[146];
	assign out[147] = registers[147];
	assign out[148] = registers[148];

	always_ff @(posedge clock) begin
		if (reset == 1) begin
			for(int i=0; i<149; i=i+1) registers[i] <= 'b0;
		end
		else begin
			registers[148:1] <= registers[147:0];
			registers[0] <= in;
		end
	end
endmodule


module counter (
	input  clock, reset,
	output logic [11:0] state,
	output logic [11:0] rev_state
);
	always_comb begin
		for (int i = 0; i < 12; i+=1) begin
			rev_state[i] = state[11-i];
		end
	end

	always_ff @(posedge clock) begin
		if (reset == 1) state <= 'b0; else
		                state <= state + 1;
	end
endmodule


module compara (
	input  logic [11:0] r,
	input  logic [11:0] p,
	output logic       out
);
	assign out = r < p;
endmodule


module compara_inv (
	input  logic [11:0] r,
	input  logic [11:0] p,
	output logic       out
);
	assign out = ~(r < p);
endmodule


module comparator_array_pos (
	input  logic [11:0] in [148:0],
	input  logic [11:0] r,
	output logic       xs [148:0]
);
	logic [11:0] r_inv;
	assign r_inv = ~r;

	compara     comp0(.r(r),     .p(in[0]), .out(xs[0]));
	compara     comp1(.r(r),     .p(in[1]), .out(xs[1]));
	compara     comp2(.r(r),     .p(in[2]), .out(xs[2]));
	compara     comp3(.r(r),     .p(in[3]), .out(xs[3]));
	compara     comp4(.r(r),     .p(in[4]), .out(xs[4]));
	compara     comp5(.r(r),     .p(in[5]), .out(xs[5]));
	compara     comp6(.r(r),     .p(in[6]), .out(xs[6]));
	compara     comp7(.r(r),     .p(in[7]), .out(xs[7]));
	compara     comp8(.r(r),     .p(in[8]), .out(xs[8]));
	compara     comp9(.r(r),     .p(in[9]), .out(xs[9]));
	compara     comp10(.r(r),     .p(in[10]), .out(xs[10]));
	compara     comp11(.r(r),     .p(in[11]), .out(xs[11]));
	compara     comp12(.r(r),     .p(in[12]), .out(xs[12]));
	compara     comp13(.r(r),     .p(in[13]), .out(xs[13]));
	compara     comp14(.r(r),     .p(in[14]), .out(xs[14]));
	compara     comp15(.r(r),     .p(in[15]), .out(xs[15]));
	compara     comp16(.r(r),     .p(in[16]), .out(xs[16]));
	compara     comp17(.r(r),     .p(in[17]), .out(xs[17]));
	compara     comp18(.r(r),     .p(in[18]), .out(xs[18]));
	compara     comp19(.r(r),     .p(in[19]), .out(xs[19]));
	compara     comp20(.r(r),     .p(in[20]), .out(xs[20]));
	compara     comp21(.r(r),     .p(in[21]), .out(xs[21]));
	compara     comp22(.r(r),     .p(in[22]), .out(xs[22]));
	compara     comp23(.r(r),     .p(in[23]), .out(xs[23]));
	compara     comp24(.r(r),     .p(in[24]), .out(xs[24]));
	compara     comp25(.r(r),     .p(in[25]), .out(xs[25]));
	compara     comp26(.r(r),     .p(in[26]), .out(xs[26]));
	compara     comp27(.r(r),     .p(in[27]), .out(xs[27]));
	compara     comp28(.r(r),     .p(in[28]), .out(xs[28]));
	compara     comp29(.r(r),     .p(in[29]), .out(xs[29]));
	compara     comp30(.r(r),     .p(in[30]), .out(xs[30]));
	compara     comp31(.r(r),     .p(in[31]), .out(xs[31]));
	compara     comp32(.r(r),     .p(in[32]), .out(xs[32]));
	compara     comp33(.r(r),     .p(in[33]), .out(xs[33]));
	compara     comp34(.r(r),     .p(in[34]), .out(xs[34]));
	compara     comp35(.r(r),     .p(in[35]), .out(xs[35]));
	compara     comp36(.r(r),     .p(in[36]), .out(xs[36]));
	compara     comp37(.r(r),     .p(in[37]), .out(xs[37]));
	compara     comp38(.r(r),     .p(in[38]), .out(xs[38]));
	compara     comp39(.r(r),     .p(in[39]), .out(xs[39]));
	compara     comp40(.r(r),     .p(in[40]), .out(xs[40]));
	compara     comp41(.r(r),     .p(in[41]), .out(xs[41]));
	compara     comp42(.r(r),     .p(in[42]), .out(xs[42]));
	compara     comp43(.r(r),     .p(in[43]), .out(xs[43]));
	compara     comp44(.r(r),     .p(in[44]), .out(xs[44]));
	compara     comp45(.r(r),     .p(in[45]), .out(xs[45]));
	compara     comp46(.r(r),     .p(in[46]), .out(xs[46]));
	compara     comp47(.r(r),     .p(in[47]), .out(xs[47]));
	compara     comp48(.r(r),     .p(in[48]), .out(xs[48]));
	compara     comp49(.r(r),     .p(in[49]), .out(xs[49]));
	compara     comp50(.r(r),     .p(in[50]), .out(xs[50]));
	compara     comp51(.r(r),     .p(in[51]), .out(xs[51]));
	compara     comp52(.r(r),     .p(in[52]), .out(xs[52]));
	compara     comp53(.r(r),     .p(in[53]), .out(xs[53]));
	compara     comp54(.r(r),     .p(in[54]), .out(xs[54]));
	compara     comp55(.r(r),     .p(in[55]), .out(xs[55]));
	compara     comp56(.r(r),     .p(in[56]), .out(xs[56]));
	compara     comp57(.r(r),     .p(in[57]), .out(xs[57]));
	compara     comp58(.r(r),     .p(in[58]), .out(xs[58]));
	compara     comp59(.r(r),     .p(in[59]), .out(xs[59]));
	compara     comp60(.r(r),     .p(in[60]), .out(xs[60]));
	compara     comp61(.r(r),     .p(in[61]), .out(xs[61]));
	compara     comp62(.r(r),     .p(in[62]), .out(xs[62]));
	compara     comp63(.r(r),     .p(in[63]), .out(xs[63]));
	compara     comp64(.r(r),     .p(in[64]), .out(xs[64]));
	compara     comp65(.r(r),     .p(in[65]), .out(xs[65]));
	compara     comp66(.r(r),     .p(in[66]), .out(xs[66]));
	compara     comp67(.r(r),     .p(in[67]), .out(xs[67]));
	compara     comp68(.r(r),     .p(in[68]), .out(xs[68]));
	compara     comp69(.r(r),     .p(in[69]), .out(xs[69]));
	compara     comp70(.r(r),     .p(in[70]), .out(xs[70]));
	compara     comp71(.r(r),     .p(in[71]), .out(xs[71]));
	compara     comp72(.r(r),     .p(in[72]), .out(xs[72]));
	compara     comp73(.r(r),     .p(in[73]), .out(xs[73]));
	compara     comp74(.r(r),     .p(in[74]), .out(xs[74]));
	compara     comp75(.r(r),     .p(in[75]), .out(xs[75]));
	compara     comp76(.r(r),     .p(in[76]), .out(xs[76]));
	compara     comp77(.r(r),     .p(in[77]), .out(xs[77]));
	compara     comp78(.r(r),     .p(in[78]), .out(xs[78]));
	compara     comp79(.r(r),     .p(in[79]), .out(xs[79]));
	compara     comp80(.r(r),     .p(in[80]), .out(xs[80]));
	compara     comp81(.r(r),     .p(in[81]), .out(xs[81]));
	compara     comp82(.r(r),     .p(in[82]), .out(xs[82]));
	compara     comp83(.r(r),     .p(in[83]), .out(xs[83]));
	compara     comp84(.r(r),     .p(in[84]), .out(xs[84]));
	compara     comp85(.r(r),     .p(in[85]), .out(xs[85]));
	compara     comp86(.r(r),     .p(in[86]), .out(xs[86]));
	compara     comp87(.r(r),     .p(in[87]), .out(xs[87]));
	compara     comp88(.r(r),     .p(in[88]), .out(xs[88]));
	compara     comp89(.r(r),     .p(in[89]), .out(xs[89]));
	compara     comp90(.r(r),     .p(in[90]), .out(xs[90]));
	compara     comp91(.r(r),     .p(in[91]), .out(xs[91]));
	compara     comp92(.r(r),     .p(in[92]), .out(xs[92]));
	compara     comp93(.r(r),     .p(in[93]), .out(xs[93]));
	compara     comp94(.r(r),     .p(in[94]), .out(xs[94]));
	compara     comp95(.r(r),     .p(in[95]), .out(xs[95]));
	compara     comp96(.r(r),     .p(in[96]), .out(xs[96]));
	compara     comp97(.r(r),     .p(in[97]), .out(xs[97]));
	compara     comp98(.r(r),     .p(in[98]), .out(xs[98]));
	compara     comp99(.r(r),     .p(in[99]), .out(xs[99]));
	compara     comp100(.r(r),     .p(in[100]), .out(xs[100]));
	compara     comp101(.r(r),     .p(in[101]), .out(xs[101]));
	compara     comp102(.r(r),     .p(in[102]), .out(xs[102]));
	compara     comp103(.r(r),     .p(in[103]), .out(xs[103]));
	compara     comp104(.r(r),     .p(in[104]), .out(xs[104]));
	compara     comp105(.r(r),     .p(in[105]), .out(xs[105]));
	compara     comp106(.r(r),     .p(in[106]), .out(xs[106]));
	compara     comp107(.r(r),     .p(in[107]), .out(xs[107]));
	compara     comp108(.r(r),     .p(in[108]), .out(xs[108]));
	compara     comp109(.r(r),     .p(in[109]), .out(xs[109]));
	compara     comp110(.r(r),     .p(in[110]), .out(xs[110]));
	compara     comp111(.r(r),     .p(in[111]), .out(xs[111]));
	compara     comp112(.r(r),     .p(in[112]), .out(xs[112]));
	compara     comp113(.r(r),     .p(in[113]), .out(xs[113]));
	compara     comp114(.r(r),     .p(in[114]), .out(xs[114]));
	compara     comp115(.r(r),     .p(in[115]), .out(xs[115]));
	compara     comp116(.r(r),     .p(in[116]), .out(xs[116]));
	compara     comp117(.r(r),     .p(in[117]), .out(xs[117]));
	compara     comp118(.r(r),     .p(in[118]), .out(xs[118]));
	compara     comp119(.r(r),     .p(in[119]), .out(xs[119]));
	compara     comp120(.r(r),     .p(in[120]), .out(xs[120]));
	compara     comp121(.r(r),     .p(in[121]), .out(xs[121]));
	compara     comp122(.r(r),     .p(in[122]), .out(xs[122]));
	compara     comp123(.r(r),     .p(in[123]), .out(xs[123]));
	compara     comp124(.r(r),     .p(in[124]), .out(xs[124]));
	compara     comp125(.r(r),     .p(in[125]), .out(xs[125]));
	compara     comp126(.r(r),     .p(in[126]), .out(xs[126]));
	compara     comp127(.r(r),     .p(in[127]), .out(xs[127]));
	compara     comp128(.r(r),     .p(in[128]), .out(xs[128]));
	compara     comp129(.r(r),     .p(in[129]), .out(xs[129]));
	compara     comp130(.r(r),     .p(in[130]), .out(xs[130]));
	compara     comp131(.r(r),     .p(in[131]), .out(xs[131]));
	compara     comp132(.r(r),     .p(in[132]), .out(xs[132]));
	compara     comp133(.r(r),     .p(in[133]), .out(xs[133]));
	compara     comp134(.r(r),     .p(in[134]), .out(xs[134]));
	compara     comp135(.r(r),     .p(in[135]), .out(xs[135]));
	compara     comp136(.r(r),     .p(in[136]), .out(xs[136]));
	compara     comp137(.r(r),     .p(in[137]), .out(xs[137]));
	compara     comp138(.r(r),     .p(in[138]), .out(xs[138]));
	compara     comp139(.r(r),     .p(in[139]), .out(xs[139]));
	compara     comp140(.r(r),     .p(in[140]), .out(xs[140]));
	compara     comp141(.r(r),     .p(in[141]), .out(xs[141]));
	compara     comp142(.r(r),     .p(in[142]), .out(xs[142]));
	compara     comp143(.r(r),     .p(in[143]), .out(xs[143]));
	compara     comp144(.r(r),     .p(in[144]), .out(xs[144]));
	compara     comp145(.r(r),     .p(in[145]), .out(xs[145]));
	compara     comp146(.r(r),     .p(in[146]), .out(xs[146]));
	compara     comp147(.r(r),     .p(in[147]), .out(xs[147]));
	compara     comp148(.r(r),     .p(in[148]), .out(xs[148]));
endmodule


module comparator_array_neg (
	input  logic [11:0] in [148:0],
	input  logic [11:0] r,
	output logic       xs [148:0]
);
	logic [11:0] r_inv;
	assign r_inv = ~r;

	compara_inv comp0(.r(r_inv), .p(in[0]), .out(xs[0]));
	compara_inv comp1(.r(r_inv), .p(in[1]), .out(xs[1]));
	compara_inv comp2(.r(r_inv), .p(in[2]), .out(xs[2]));
	compara_inv comp3(.r(r_inv), .p(in[3]), .out(xs[3]));
	compara_inv comp4(.r(r_inv), .p(in[4]), .out(xs[4]));
	compara_inv comp5(.r(r_inv), .p(in[5]), .out(xs[5]));
	compara_inv comp6(.r(r_inv), .p(in[6]), .out(xs[6]));
	compara_inv comp7(.r(r_inv), .p(in[7]), .out(xs[7]));
	compara_inv comp8(.r(r_inv), .p(in[8]), .out(xs[8]));
	compara_inv comp9(.r(r_inv), .p(in[9]), .out(xs[9]));
	compara_inv comp10(.r(r_inv), .p(in[10]), .out(xs[10]));
	compara_inv comp11(.r(r_inv), .p(in[11]), .out(xs[11]));
	compara_inv comp12(.r(r_inv), .p(in[12]), .out(xs[12]));
	compara_inv comp13(.r(r_inv), .p(in[13]), .out(xs[13]));
	compara_inv comp14(.r(r_inv), .p(in[14]), .out(xs[14]));
	compara_inv comp15(.r(r_inv), .p(in[15]), .out(xs[15]));
	compara_inv comp16(.r(r_inv), .p(in[16]), .out(xs[16]));
	compara_inv comp17(.r(r_inv), .p(in[17]), .out(xs[17]));
	compara_inv comp18(.r(r_inv), .p(in[18]), .out(xs[18]));
	compara_inv comp19(.r(r_inv), .p(in[19]), .out(xs[19]));
	compara_inv comp20(.r(r_inv), .p(in[20]), .out(xs[20]));
	compara_inv comp21(.r(r_inv), .p(in[21]), .out(xs[21]));
	compara_inv comp22(.r(r_inv), .p(in[22]), .out(xs[22]));
	compara_inv comp23(.r(r_inv), .p(in[23]), .out(xs[23]));
	compara_inv comp24(.r(r_inv), .p(in[24]), .out(xs[24]));
	compara_inv comp25(.r(r_inv), .p(in[25]), .out(xs[25]));
	compara_inv comp26(.r(r_inv), .p(in[26]), .out(xs[26]));
	compara_inv comp27(.r(r_inv), .p(in[27]), .out(xs[27]));
	compara_inv comp28(.r(r_inv), .p(in[28]), .out(xs[28]));
	compara_inv comp29(.r(r_inv), .p(in[29]), .out(xs[29]));
	compara_inv comp30(.r(r_inv), .p(in[30]), .out(xs[30]));
	compara_inv comp31(.r(r_inv), .p(in[31]), .out(xs[31]));
	compara_inv comp32(.r(r_inv), .p(in[32]), .out(xs[32]));
	compara_inv comp33(.r(r_inv), .p(in[33]), .out(xs[33]));
	compara_inv comp34(.r(r_inv), .p(in[34]), .out(xs[34]));
	compara_inv comp35(.r(r_inv), .p(in[35]), .out(xs[35]));
	compara_inv comp36(.r(r_inv), .p(in[36]), .out(xs[36]));
	compara_inv comp37(.r(r_inv), .p(in[37]), .out(xs[37]));
	compara_inv comp38(.r(r_inv), .p(in[38]), .out(xs[38]));
	compara_inv comp39(.r(r_inv), .p(in[39]), .out(xs[39]));
	compara_inv comp40(.r(r_inv), .p(in[40]), .out(xs[40]));
	compara_inv comp41(.r(r_inv), .p(in[41]), .out(xs[41]));
	compara_inv comp42(.r(r_inv), .p(in[42]), .out(xs[42]));
	compara_inv comp43(.r(r_inv), .p(in[43]), .out(xs[43]));
	compara_inv comp44(.r(r_inv), .p(in[44]), .out(xs[44]));
	compara_inv comp45(.r(r_inv), .p(in[45]), .out(xs[45]));
	compara_inv comp46(.r(r_inv), .p(in[46]), .out(xs[46]));
	compara_inv comp47(.r(r_inv), .p(in[47]), .out(xs[47]));
	compara_inv comp48(.r(r_inv), .p(in[48]), .out(xs[48]));
	compara_inv comp49(.r(r_inv), .p(in[49]), .out(xs[49]));
	compara_inv comp50(.r(r_inv), .p(in[50]), .out(xs[50]));
	compara_inv comp51(.r(r_inv), .p(in[51]), .out(xs[51]));
	compara_inv comp52(.r(r_inv), .p(in[52]), .out(xs[52]));
	compara_inv comp53(.r(r_inv), .p(in[53]), .out(xs[53]));
	compara_inv comp54(.r(r_inv), .p(in[54]), .out(xs[54]));
	compara_inv comp55(.r(r_inv), .p(in[55]), .out(xs[55]));
	compara_inv comp56(.r(r_inv), .p(in[56]), .out(xs[56]));
	compara_inv comp57(.r(r_inv), .p(in[57]), .out(xs[57]));
	compara_inv comp58(.r(r_inv), .p(in[58]), .out(xs[58]));
	compara_inv comp59(.r(r_inv), .p(in[59]), .out(xs[59]));
	compara_inv comp60(.r(r_inv), .p(in[60]), .out(xs[60]));
	compara_inv comp61(.r(r_inv), .p(in[61]), .out(xs[61]));
	compara_inv comp62(.r(r_inv), .p(in[62]), .out(xs[62]));
	compara_inv comp63(.r(r_inv), .p(in[63]), .out(xs[63]));
	compara_inv comp64(.r(r_inv), .p(in[64]), .out(xs[64]));
	compara_inv comp65(.r(r_inv), .p(in[65]), .out(xs[65]));
	compara_inv comp66(.r(r_inv), .p(in[66]), .out(xs[66]));
	compara_inv comp67(.r(r_inv), .p(in[67]), .out(xs[67]));
	compara_inv comp68(.r(r_inv), .p(in[68]), .out(xs[68]));
	compara_inv comp69(.r(r_inv), .p(in[69]), .out(xs[69]));
	compara_inv comp70(.r(r_inv), .p(in[70]), .out(xs[70]));
	compara_inv comp71(.r(r_inv), .p(in[71]), .out(xs[71]));
	compara_inv comp72(.r(r_inv), .p(in[72]), .out(xs[72]));
	compara_inv comp73(.r(r_inv), .p(in[73]), .out(xs[73]));
	compara_inv comp74(.r(r_inv), .p(in[74]), .out(xs[74]));
	compara_inv comp75(.r(r_inv), .p(in[75]), .out(xs[75]));
	compara_inv comp76(.r(r_inv), .p(in[76]), .out(xs[76]));
	compara_inv comp77(.r(r_inv), .p(in[77]), .out(xs[77]));
	compara_inv comp78(.r(r_inv), .p(in[78]), .out(xs[78]));
	compara_inv comp79(.r(r_inv), .p(in[79]), .out(xs[79]));
	compara_inv comp80(.r(r_inv), .p(in[80]), .out(xs[80]));
	compara_inv comp81(.r(r_inv), .p(in[81]), .out(xs[81]));
	compara_inv comp82(.r(r_inv), .p(in[82]), .out(xs[82]));
	compara_inv comp83(.r(r_inv), .p(in[83]), .out(xs[83]));
	compara_inv comp84(.r(r_inv), .p(in[84]), .out(xs[84]));
	compara_inv comp85(.r(r_inv), .p(in[85]), .out(xs[85]));
	compara_inv comp86(.r(r_inv), .p(in[86]), .out(xs[86]));
	compara_inv comp87(.r(r_inv), .p(in[87]), .out(xs[87]));
	compara_inv comp88(.r(r_inv), .p(in[88]), .out(xs[88]));
	compara_inv comp89(.r(r_inv), .p(in[89]), .out(xs[89]));
	compara_inv comp90(.r(r_inv), .p(in[90]), .out(xs[90]));
	compara_inv comp91(.r(r_inv), .p(in[91]), .out(xs[91]));
	compara_inv comp92(.r(r_inv), .p(in[92]), .out(xs[92]));
	compara_inv comp93(.r(r_inv), .p(in[93]), .out(xs[93]));
	compara_inv comp94(.r(r_inv), .p(in[94]), .out(xs[94]));
	compara_inv comp95(.r(r_inv), .p(in[95]), .out(xs[95]));
	compara_inv comp96(.r(r_inv), .p(in[96]), .out(xs[96]));
	compara_inv comp97(.r(r_inv), .p(in[97]), .out(xs[97]));
	compara_inv comp98(.r(r_inv), .p(in[98]), .out(xs[98]));
	compara_inv comp99(.r(r_inv), .p(in[99]), .out(xs[99]));
	compara_inv comp100(.r(r_inv), .p(in[100]), .out(xs[100]));
	compara_inv comp101(.r(r_inv), .p(in[101]), .out(xs[101]));
	compara_inv comp102(.r(r_inv), .p(in[102]), .out(xs[102]));
	compara_inv comp103(.r(r_inv), .p(in[103]), .out(xs[103]));
	compara_inv comp104(.r(r_inv), .p(in[104]), .out(xs[104]));
	compara_inv comp105(.r(r_inv), .p(in[105]), .out(xs[105]));
	compara_inv comp106(.r(r_inv), .p(in[106]), .out(xs[106]));
	compara_inv comp107(.r(r_inv), .p(in[107]), .out(xs[107]));
	compara_inv comp108(.r(r_inv), .p(in[108]), .out(xs[108]));
	compara_inv comp109(.r(r_inv), .p(in[109]), .out(xs[109]));
	compara_inv comp110(.r(r_inv), .p(in[110]), .out(xs[110]));
	compara_inv comp111(.r(r_inv), .p(in[111]), .out(xs[111]));
	compara_inv comp112(.r(r_inv), .p(in[112]), .out(xs[112]));
	compara_inv comp113(.r(r_inv), .p(in[113]), .out(xs[113]));
	compara_inv comp114(.r(r_inv), .p(in[114]), .out(xs[114]));
	compara_inv comp115(.r(r_inv), .p(in[115]), .out(xs[115]));
	compara_inv comp116(.r(r_inv), .p(in[116]), .out(xs[116]));
	compara_inv comp117(.r(r_inv), .p(in[117]), .out(xs[117]));
	compara_inv comp118(.r(r_inv), .p(in[118]), .out(xs[118]));
	compara_inv comp119(.r(r_inv), .p(in[119]), .out(xs[119]));
	compara_inv comp120(.r(r_inv), .p(in[120]), .out(xs[120]));
	compara_inv comp121(.r(r_inv), .p(in[121]), .out(xs[121]));
	compara_inv comp122(.r(r_inv), .p(in[122]), .out(xs[122]));
	compara_inv comp123(.r(r_inv), .p(in[123]), .out(xs[123]));
	compara_inv comp124(.r(r_inv), .p(in[124]), .out(xs[124]));
	compara_inv comp125(.r(r_inv), .p(in[125]), .out(xs[125]));
	compara_inv comp126(.r(r_inv), .p(in[126]), .out(xs[126]));
	compara_inv comp127(.r(r_inv), .p(in[127]), .out(xs[127]));
	compara_inv comp128(.r(r_inv), .p(in[128]), .out(xs[128]));
	compara_inv comp129(.r(r_inv), .p(in[129]), .out(xs[129]));
	compara_inv comp130(.r(r_inv), .p(in[130]), .out(xs[130]));
	compara_inv comp131(.r(r_inv), .p(in[131]), .out(xs[131]));
	compara_inv comp132(.r(r_inv), .p(in[132]), .out(xs[132]));
	compara_inv comp133(.r(r_inv), .p(in[133]), .out(xs[133]));
	compara_inv comp134(.r(r_inv), .p(in[134]), .out(xs[134]));
	compara_inv comp135(.r(r_inv), .p(in[135]), .out(xs[135]));
	compara_inv comp136(.r(r_inv), .p(in[136]), .out(xs[136]));
	compara_inv comp137(.r(r_inv), .p(in[137]), .out(xs[137]));
	compara_inv comp138(.r(r_inv), .p(in[138]), .out(xs[138]));
	compara_inv comp139(.r(r_inv), .p(in[139]), .out(xs[139]));
	compara_inv comp140(.r(r_inv), .p(in[140]), .out(xs[140]));
	compara_inv comp141(.r(r_inv), .p(in[141]), .out(xs[141]));
	compara_inv comp142(.r(r_inv), .p(in[142]), .out(xs[142]));
	compara_inv comp143(.r(r_inv), .p(in[143]), .out(xs[143]));
	compara_inv comp144(.r(r_inv), .p(in[144]), .out(xs[144]));
	compara_inv comp145(.r(r_inv), .p(in[145]), .out(xs[145]));
	compara_inv comp146(.r(r_inv), .p(in[146]), .out(xs[146]));
	compara_inv comp147(.r(r_inv), .p(in[147]), .out(xs[147]));
	compara_inv comp148(.r(r_inv), .p(in[148]), .out(xs[148]));
endmodule


module hw_tree0  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[2] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[3] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[4] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[5] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[6] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[7] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[8] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[9] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[10] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[11] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[12] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[13] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[14] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[15] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[16] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[17] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[18] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[19] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[20] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[21] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[22] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[23] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[24] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[25] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[26] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[27] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[28] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[29] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[30] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[31] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[32] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[33] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[34] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[35] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[36] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[37] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[38] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[39] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[40] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[41] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[42] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[43] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[44] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[45] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[46] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[47] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[48] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[49] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[50] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[51] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[52] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[53] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[54] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[55] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[56] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[57] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[58] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[59] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[60] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[61] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[62] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[63] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[64] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[65] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[66] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[67] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[68] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[69] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[70] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[71] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[72] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[73] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[74] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[75] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[76] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[77] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[78] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[79] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[80] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[81] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[82] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[83] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[84] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[85] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[86] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[87] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[88] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[89] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[90] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[91] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[92] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[93] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[94] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[95] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[96] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[97] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[98] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[99] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[100] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[101] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[102] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[103] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[104] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[105] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[106] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[107] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[108] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[109] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[110] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[111] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[112] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[113] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[114] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[115] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[116] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[117] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[118] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[119] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[120] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[121] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[122] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[123] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[124] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[125] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[126] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[127] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[128] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[129] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[130] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[131] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[132] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[133] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[134] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[135] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[136] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[137] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[138] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[139] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[140] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[141] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[142] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[143] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[144] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[145] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[146] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[147] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[148] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[149] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[150] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[151] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[152] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[153] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[154] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[155] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[156] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[157] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[158] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[159] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[160] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[161] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[162] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[163] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[164] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[165] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[166] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[167] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[168] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[169] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[170] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[171] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[172] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[173] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[174] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[175] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[176] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[177] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[178] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[179] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[180] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[181] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[182] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[183] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[184] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[185] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[186] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[187] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[188] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[189] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[190] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[191] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[192] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[193] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[194] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[195] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[196] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[197] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[198] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[199] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[200] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[201] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[202] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[203] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[204] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[205] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[206] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[207] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[208] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[209] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[210] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[211] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[212] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[213] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[214] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[215] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[216] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[217] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[218] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[219] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[220] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[221] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[222] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[223] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[224] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[225] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[226] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[227] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[228] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[229] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[230] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[231] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[232] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[233] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[234] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[235] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[236] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[237] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[238] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[239] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[240] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[241] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[242] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[243] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[244] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[245] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[246] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[247] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[248] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[249] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[250] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[251] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[252] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[253] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[254] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[255] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[256] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[257] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[258] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[259] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[260] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[261] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[262] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[263] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[264] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[265] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[266] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[267] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[268] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[269] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[270] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[271] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[272] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[273] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[274] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[275] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[276] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[277] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[278] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[279] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[280] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[281] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[282] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[283] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[284] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[285] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[286] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[287] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[288] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[289] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[290] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[291] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[292] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[293] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[294] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[295] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[296] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[297] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[298] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[299] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[300] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[301] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[302] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[303] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[304] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[305] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[306] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[307] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[308] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[309] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[310] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[311] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[312] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[313] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[314] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[315] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[316] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[317] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[318] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[319] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[320] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[321] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[322] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[323] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[324] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[325] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[326] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[327] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[328] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[329] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[330] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[331] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[332] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[333] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[334] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[335] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[336] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[337] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[338] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[339] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[340] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[341] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[342] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[343] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[344] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[345] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[346] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[347] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[348] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[349] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[350] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[351] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[352] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[353] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[354] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[355] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[356] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[357] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[358] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[359] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[360] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[361] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[362] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[363] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[364] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[365] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[366] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[367] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[368] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[369] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[370] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[371] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[372] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[373] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[374] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[375] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[376] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[377] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[378] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[379] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[380] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[381] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[382] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[383] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[384] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[385] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[386] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[387] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[388] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[389] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[390] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[391] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[392] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[393] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[394] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[395] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[396] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[397] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[398] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[399] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[400] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[401] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[402] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[403] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[404] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[405] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[406] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[407] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[408] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[409] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[410] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[411] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[412] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[413] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[414] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[415] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[416] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[417] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[418] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[419] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[420] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[421] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[422] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[423] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[424] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[425] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[426] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[427] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[428] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[429] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[430] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[431] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[432] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[433] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[434] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[435] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[436] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[437] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[438] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[439] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[440] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[441] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[442] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[443] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[444] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[445] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[446] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[447] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[448] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[449] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[450] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[451] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[452] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[453] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[454] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[455] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[456] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[457] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[458] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[459] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[460] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[461] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[462] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[463] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[464] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[465] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[466] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[467] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[468] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[469] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[470] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[471] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[472] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[473] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[474] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[475] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[476] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[477] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[478] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[479] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[480] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[481] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[482] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[483] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[484] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[485] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[486] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[487] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[488] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[489] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[490] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[491] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[492] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[493] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[494] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[495] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[496] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[497] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[498] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[499] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[500] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[501] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[502] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[503] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[504] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[505] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[506] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[507] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[508] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[509] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[510] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[511] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[512] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[513] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[514] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[515] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[516] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[517] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[518] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[519] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[520] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[521] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[522] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[523] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[524] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[525] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[526] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[527] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[528] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[529] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[530] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[531] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[532] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[533] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[534] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[535] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[536] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[537] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[538] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[539] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[540] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[541] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[542] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[543] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[544] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[545] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[546] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[547] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[548] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[549] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[550] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[551] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[552] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[553] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[554] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[555] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[556] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[557] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[558] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[559] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[560] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[561] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[562] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[563] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[564] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[565] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[566] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[567] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[568] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[569] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[570] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[571] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[572] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[573] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[574] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[575] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[576] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[577] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[578] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[579] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[580] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[581] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[582] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[583] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[584] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[585] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[586] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[587] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[588] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[589] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[590] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[591] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[592] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[593] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[594] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[595] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[596] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[597] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[598] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[599] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[600] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[601] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[602] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[603] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[604] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[605] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[606] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[607] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[608] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[609] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[610] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[611] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[612] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[613] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[614] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[615] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[616] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[617] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[618] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[619] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[620] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[621] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[622] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[623] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[624] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[625] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[626] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[627] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[628] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[629] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[630] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[631] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[632] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[633] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[634] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[635] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[636] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[637] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[638] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[639] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[640] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[641] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[642] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[643] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[644] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[645] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[646] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[647] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[648] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[649] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[650] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[651] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[652] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[653] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[654] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[655] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[656] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[657] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[658] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[659] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[660] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[661] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[662] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[663] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[664] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[665] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[666] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[667] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[668] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[669] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[670] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[671] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[672] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[673] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[674] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[675] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[676] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[677] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[678] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[679] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[680] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[681] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[682] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[683] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[684] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[685] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[686] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[687] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[688] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[689] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[690] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[691] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[692] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[693] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[694] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[695] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[696] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[697] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[698] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[699] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[700] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[701] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[702] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[703] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[704] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[705] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[706] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[707] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[708] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[709] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[710] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[711] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[712] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[713] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[714] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[715] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[716] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[717] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[718] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[719] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[720] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[721] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[722] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[723] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[724] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[725] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[726] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[727] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[728] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[729] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[730] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[731] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[732] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[733] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[734] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[735] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[736] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[737] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[738] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[739] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[740] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[741] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[742] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[743] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[744] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[745] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[746] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[747] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[748] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[749] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[750] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[751] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[752] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[753] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[754] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[755] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[756] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[757] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[758] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[759] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[760] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[761] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[762] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[763] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[764] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[765] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[766] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[767] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[768] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[769] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[770] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[771] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[772] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[773] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[774] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[775] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[776] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[777] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[778] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[779] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[780] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[781] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[782] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[783] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[784] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[785] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[786] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[787] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[788] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[789] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[790] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[791] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[792] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[793] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[794] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[795] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[796] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[797] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[798] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[799] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[800] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[801] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[802] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[803] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[804] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[805] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[806] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[807] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[808] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[809] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[810] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[811] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[812] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[813] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[814] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[815] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[816] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[817] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[818] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[819] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[820] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[821] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[822] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[823] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[824] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[825] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[826] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[827] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[828] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[829] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[830] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[831] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[832] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[833] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[834] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[835] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[836] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[837] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[838] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[839] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[840] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[841] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[842] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[843] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[844] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[845] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[846] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[847] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[848] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[849] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[850] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[851] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[852] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[853] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[854] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[855] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[856] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[857] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[858] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[859] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[860] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[861] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[862] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[863] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[864] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[865] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[866] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[867] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[868] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[869] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[870] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[871] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[872] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[873] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[874] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[875] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[876] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[877] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[878] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[879] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[880] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[881] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[882] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[883] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[884] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[885] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[886] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[887] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[888] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[889] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[890] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[891] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[892] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[893] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[894] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[895] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[896] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[897] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[898] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[899] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[900] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[901] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[902] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[903] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[904] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[905] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[906] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[907] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[908] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[909] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[910] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[911] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[912] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[913] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[914] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[915] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[916] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[917] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[918] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[919] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[920] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[921] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[922] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[923] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[924] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[925] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[926] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[927] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[928] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[929] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[930] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[931] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[932] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[933] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[934] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[935] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[936] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[937] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[938] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[939] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[940] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[941] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[942] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[943] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[944] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[945] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[946] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[947] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[948] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[949] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[950] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[951] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[952] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[953] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[954] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[955] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[956] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[957] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[958] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[959] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[960] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[961] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[962] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[963] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[964] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[965] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[966] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[967] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[968] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[969] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[970] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[971] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[972] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[973] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[974] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[975] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[976] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[977] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[978] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[979] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[980] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[981] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[982] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[983] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[984] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[985] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[986] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[987] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[988] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[989] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[990] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[991] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[992] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[993] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[994] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[995] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[996] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[997] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[998] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[999] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1000] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1001] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1002] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1003] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1004] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1005] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1006] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1007] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1008] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1009] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1010] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1011] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1012] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1013] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1014] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1015] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1016] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1017] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1018] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1019] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1020] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1021] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1022] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1023] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1024] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1025] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1026] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1027] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1028] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1029] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1030] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1031] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1032] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1033] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1034] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1035] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1036] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1037] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1038] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1039] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1040] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1041] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1042] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1043] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1044] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1045] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1046] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1047] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1048] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1049] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1050] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1051] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1052] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1053] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1054] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1055] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1056] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1057] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1058] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1059] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1060] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1061] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1062] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1063] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1064] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1065] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1066] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1067] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1068] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1069] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1070] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1071] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1072] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1073] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1074] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1075] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1076] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1077] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1078] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1079] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1080] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1081] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1082] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1083] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1084] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1085] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1086] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1087] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1088] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1089] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1090] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1091] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1092] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1093] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1094] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1095] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1096] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1097] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1098] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1099] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1100] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1101] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1102] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1103] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1104] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1105] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1106] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1107] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1108] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1109] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1110] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1111] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1112] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1113] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1114] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1115] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1116] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1117] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1118] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1119] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1120] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1121] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1122] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1123] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1124] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1125] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1126] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1127] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1128] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1129] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1130] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1131] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1132] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1133] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1134] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1135] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1136] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1137] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1138] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1139] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1140] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1141] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1142] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1143] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1144] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1145] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1146] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1147] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1148] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1149] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1150] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1151] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1152] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1153] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1154] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1155] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1156] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1157] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1158] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1159] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1160] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1161] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1162] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1163] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1164] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1165] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1166] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1167] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1168] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1169] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1170] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1171] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1172] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1173] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1174] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1175] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1176] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1177] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1178] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1179] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1180] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1181] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1182] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1183] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1184] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1185] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1186] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1187] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1188] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1189] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1190] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1191] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1192] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1193] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1194] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1195] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1196] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1197] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1198] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1199] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1200] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1201] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1202] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1203] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1204] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1205] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1206] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1207] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1208] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1209] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1210] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1211] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1212] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1213] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1214] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1215] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1216] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1217] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1218] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1219] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1220] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1221] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1222] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1223] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1224] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1225] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1226] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1227] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1228] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1229] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1230] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1231] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1232] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1233] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1234] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1235] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1236] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1237] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1238] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1239] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1240] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1241] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1242] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1243] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1244] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1245] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1246] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1247] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1248] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1249] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1250] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1251] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1252] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1253] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1254] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1255] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1256] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1257] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1258] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1259] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1260] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1261] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1262] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1263] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1264] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1265] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1266] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1267] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1268] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1269] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1270] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1271] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1272] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1273] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1274] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1275] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1276] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1277] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1278] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1279] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1280] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1281] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1282] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1283] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1284] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1285] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1286] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1287] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1288] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1289] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1290] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1291] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1292] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1293] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1294] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1295] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1296] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1297] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1298] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1299] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1300] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1301] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1302] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1303] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1304] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1305] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1306] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1307] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1308] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1309] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1310] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1311] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1312] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1313] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1314] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1315] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1316] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1317] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1318] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1319] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1320] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1321] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1322] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1323] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1324] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1325] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1326] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1327] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1328] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1329] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1330] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1331] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1332] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1333] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1334] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1335] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1336] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1337] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1338] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1339] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1340] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1341] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1342] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1343] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1344] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1345] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1346] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1347] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1348] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1349] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1350] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1351] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1352] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1353] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1354] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1355] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1356] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1357] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1358] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1359] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1360] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1361] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1362] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1363] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1364] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1365] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1366] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1367] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1368] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1369] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1370] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1371] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1372] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1373] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1374] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1375] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1376] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1377] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1378] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1379] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1380] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1381] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1382] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1383] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1384] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1385] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1386] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1387] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1388] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1389] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1390] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1391] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1392] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1393] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1394] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1395] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1396] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1397] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1398] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1399] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1400] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1401] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1402] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1403] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1404] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1405] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1406] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1407] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1408] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1409] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1410] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1411] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1412] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1413] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1414] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1415] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1416] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1417] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1418] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1419] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1420] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1421] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1422] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1423] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1424] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1425] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1426] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1427] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1428] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1429] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1430] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1431] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1432] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1433] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1434] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1435] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1436] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1437] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1438] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1439] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1440] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1441] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1442] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1443] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1444] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1445] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1446] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1447] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1448] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1449] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1450] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1451] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1452] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1453] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1454] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1455] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1456] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1457] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1458] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1459] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1460] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1461] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1462] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1463] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1464] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1465] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1466] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1467] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1468] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1469] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1470] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1471] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1472] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1473] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1474] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1475] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1476] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1477] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1478] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1479] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1480] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1481] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1482] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1483] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1484] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1485] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1486] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1487] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1488] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1489] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1490] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1491] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1492] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1493] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1494] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1495] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1496] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1497] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1498] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1499] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1500] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1501] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1502] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1503] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1504] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1505] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1506] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1507] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1508] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1509] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1510] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1511] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1512] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1513] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1514] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1515] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1516] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1517] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1518] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1519] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1520] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1521] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1522] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1523] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1524] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1525] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1526] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1527] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1528] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1529] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1530] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1531] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1532] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1533] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1534] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1535] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1536] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1537] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1538] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1539] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1540] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1541] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1542] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1543] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1544] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1545] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1546] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1547] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1548] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1549] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1550] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1551] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1552] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1553] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1554] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1555] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1556] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1557] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1558] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1559] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1560] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1561] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1562] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1563] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1564] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1565] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1566] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1567] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1568] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1569] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1570] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1571] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1572] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1573] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1574] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1575] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1576] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1577] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1578] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1579] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1580] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1581] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1582] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1583] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1584] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1585] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1586] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1587] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1588] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1589] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1590] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1591] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1592] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1593] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1594] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1595] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1596] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1597] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1598] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1599] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1600] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1601] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1602] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1603] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1604] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1605] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1606] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1607] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1608] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1609] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1610] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1611] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1612] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1613] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1614] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1615] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1616] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1617] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1618] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1619] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1620] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1621] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1622] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1623] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1624] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1625] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1626] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1627] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1628] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1629] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1630] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1631] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1632] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1633] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1634] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1635] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1636] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1637] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1638] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1639] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1640] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1641] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1642] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1643] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1644] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1645] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1646] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1647] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1648] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1649] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1650] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1651] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1652] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1653] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1654] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1655] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1656] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1657] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1658] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1659] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1660] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1661] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1662] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1663] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1664] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1665] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1666] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1667] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1668] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1669] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1670] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1671] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1672] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1673] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1674] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1675] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1676] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1677] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1678] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1679] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1680] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1681] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1682] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1683] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1684] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1685] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1686] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1687] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1688] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1689] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1690] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1691] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1692] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1693] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1694] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1695] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1696] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[1697] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[1698] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[1699] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[1700] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1701] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1702] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1703] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1704] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[1705] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[1706] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[1707] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[1708] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1709] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1710] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1711] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1712] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1713] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1714] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1715] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1716] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1717] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1718] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1719] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1720] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1721] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1722] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1723] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1724] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1725] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1726] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1727] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1728] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1729] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1730] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1731] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1732] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1733] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1734] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1735] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1736] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1737] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1738] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1739] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1740] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1741] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1742] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1743] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1744] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1745] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1746] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1747] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1748] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1749] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1750] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1751] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1752] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1753] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1754] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1755] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1756] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1757] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1758] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1759] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1760] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1761] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1762] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1763] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1764] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1765] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1766] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1767] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1768] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1769] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1770] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1771] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1772] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1773] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1774] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1775] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1776] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1777] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1778] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1779] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1780] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1781] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1782] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1783] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1784] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1785] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1786] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1787] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1788] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1789] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1790] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1791] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1792] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1793] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1794] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1795] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1796] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1797] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1798] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1799] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1800] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1801] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1802] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1803] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1804] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1805] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1806] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1807] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1808] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1809] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1810] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1811] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1812] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1813] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1814] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1815] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1816] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1817] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1818] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1819] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1820] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1821] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1822] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1823] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1824] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1825] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1826] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1827] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1828] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1829] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1830] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1831] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1832] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1833] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1834] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1835] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1836] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1837] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1838] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1839] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1840] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1841] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1842] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1843] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1844] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1845] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1846] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1847] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1848] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1849] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1850] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1851] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1852] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1853] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1854] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1855] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1856] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1857] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1858] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1859] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1860] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1861] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1862] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1863] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1864] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1865] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1866] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1867] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1868] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1869] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1870] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1871] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1872] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[1873] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[1874] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[1875] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[1876] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1877] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1878] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1879] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1880] = s[0] ? pos_SNs[111] : pos_SNs[111];
	assign level0[1881] = s[0] ? pos_SNs[111] : pos_SNs[111];
	assign level0[1882] = s[0] ? pos_SNs[111] : pos_SNs[111];
	assign level0[1883] = s[0] ? pos_SNs[111] : pos_SNs[111];
	assign level0[1884] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1885] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1886] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1887] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1888] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1889] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1890] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1891] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1892] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1893] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1894] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1895] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1896] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1897] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1898] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1899] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1900] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1901] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1902] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1903] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1904] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1905] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1906] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1907] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1908] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1909] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1910] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1911] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1912] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1913] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1914] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1915] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1916] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1917] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1918] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1919] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1920] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1921] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1922] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1923] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1924] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1925] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1926] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1927] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1928] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1929] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1930] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1931] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1932] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1933] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1934] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1935] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1936] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1937] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1938] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1939] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1940] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1941] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1942] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1943] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1944] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1945] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1946] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1947] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1948] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1949] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1950] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1951] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1952] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1953] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1954] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1955] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1956] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1957] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1958] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1959] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1960] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1961] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1962] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1963] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1964] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1965] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1966] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1967] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1968] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1969] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1970] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1971] = s[0] ? neg_SNs[28] : neg_SNs[28];
	assign level0[1972] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1973] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1974] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1975] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1976] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[1977] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1978] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1979] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1980] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1981] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1982] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1983] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1984] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1985] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1986] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1987] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1988] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1989] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1990] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1991] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1992] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1993] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1994] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1995] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1996] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1997] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1998] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1999] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[2000] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[2001] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[2002] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[2003] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[2004] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[2005] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[2006] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[2007] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[2008] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[2009] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[2010] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[2011] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[2012] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[2013] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[2014] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[2015] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2016] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[2017] = s[0] ? neg_SNs[12] : neg_SNs[12];
	assign level0[2018] = s[0] ? neg_SNs[14] : neg_SNs[14];
	assign level0[2019] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[2020] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[2021] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[2022] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[2023] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[2024] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[2025] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[2026] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[2027] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[2028] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[2029] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[2030] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[2031] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[2032] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[2033] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[2034] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[2035] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[2036] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[2037] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[2038] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[2039] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[2040] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[2041] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[2042] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[2043] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[2044] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2045] = s[0] ? neg_SNs[131] : neg_SNs[131];
	assign level0[2046] = s[0] ? neg_SNs[133] : neg_SNs[133];
	assign level0[2047] = s[0] ? neg_SNs[135] : neg_SNs[135];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module hw_tree1  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[2] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[3] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[4] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[5] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[6] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[7] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[8] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[9] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[10] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[11] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[12] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[13] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[14] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[15] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[16] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[17] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[18] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[19] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[20] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[21] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[22] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[23] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[24] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[25] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[26] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[27] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[28] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[29] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[30] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[31] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[32] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[33] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[34] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[35] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[36] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[37] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[38] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[39] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[40] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[41] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[42] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[43] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[44] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[45] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[46] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[47] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[48] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[49] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[50] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[51] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[52] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[53] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[54] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[55] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[56] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[57] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[58] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[59] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[60] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[61] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[62] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[63] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[64] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[65] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[66] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[67] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[68] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[69] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[70] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[71] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[72] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[73] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[74] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[75] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[76] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[77] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[78] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[79] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[80] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[81] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[82] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[83] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[84] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[85] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[86] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[87] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[88] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[89] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[90] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[91] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[92] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[93] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[94] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[95] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[96] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[97] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[98] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[99] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[100] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[101] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[102] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[103] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[104] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[105] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[106] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[107] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[108] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[109] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[110] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[111] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[112] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[113] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[114] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[115] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[116] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[117] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[118] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[119] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[120] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[121] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[122] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[123] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[124] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[125] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[126] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[127] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[128] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[129] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[130] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[131] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[132] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[133] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[134] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[135] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[136] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[137] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[138] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[139] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[140] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[141] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[142] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[143] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[144] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[145] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[146] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[147] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[148] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[149] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[150] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[151] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[152] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[153] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[154] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[155] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[156] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[157] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[158] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[159] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[160] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[161] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[162] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[163] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[164] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[165] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[166] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[167] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[168] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[169] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[170] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[171] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[172] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[173] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[174] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[175] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[176] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[177] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[178] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[179] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[180] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[181] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[182] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[183] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[184] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[185] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[186] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[187] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[188] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[189] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[190] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[191] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[192] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[193] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[194] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[195] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[196] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[197] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[198] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[199] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[200] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[201] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[202] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[203] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[204] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[205] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[206] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[207] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[208] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[209] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[210] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[211] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[212] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[213] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[214] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[215] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[216] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[217] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[218] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[219] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[220] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[221] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[222] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[223] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[224] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[225] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[226] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[227] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[228] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[229] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[230] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[231] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[232] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[233] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[234] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[235] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[236] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[237] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[238] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[239] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[240] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[241] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[242] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[243] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[244] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[245] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[246] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[247] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[248] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[249] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[250] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[251] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[252] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[253] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[254] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[255] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[256] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[257] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[258] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[259] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[260] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[261] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[262] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[263] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[264] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[265] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[266] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[267] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[268] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[269] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[270] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[271] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[272] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[273] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[274] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[275] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[276] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[277] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[278] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[279] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[280] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[281] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[282] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[283] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[284] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[285] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[286] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[287] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[288] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[289] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[290] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[291] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[292] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[293] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[294] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[295] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[296] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[297] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[298] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[299] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[300] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[301] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[302] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[303] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[304] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[305] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[306] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[307] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[308] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[309] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[310] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[311] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[312] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[313] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[314] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[315] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[316] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[317] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[318] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[319] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[320] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[321] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[322] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[323] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[324] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[325] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[326] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[327] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[328] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[329] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[330] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[331] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[332] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[333] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[334] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[335] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[336] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[337] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[338] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[339] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[340] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[341] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[342] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[343] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[344] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[345] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[346] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[347] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[348] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[349] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[350] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[351] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[352] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[353] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[354] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[355] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[356] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[357] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[358] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[359] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[360] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[361] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[362] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[363] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[364] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[365] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[366] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[367] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[368] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[369] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[370] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[371] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[372] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[373] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[374] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[375] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[376] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[377] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[378] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[379] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[380] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[381] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[382] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[383] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[384] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[385] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[386] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[387] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[388] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[389] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[390] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[391] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[392] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[393] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[394] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[395] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[396] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[397] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[398] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[399] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[400] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[401] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[402] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[403] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[404] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[405] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[406] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[407] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[408] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[409] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[410] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[411] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[412] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[413] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[414] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[415] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[416] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[417] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[418] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[419] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[420] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[421] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[422] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[423] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[424] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[425] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[426] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[427] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[428] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[429] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[430] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[431] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[432] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[433] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[434] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[435] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[436] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[437] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[438] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[439] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[440] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[441] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[442] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[443] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[444] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[445] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[446] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[447] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[448] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[449] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[450] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[451] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[452] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[453] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[454] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[455] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[456] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[457] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[458] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[459] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[460] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[461] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[462] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[463] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[464] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[465] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[466] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[467] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[468] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[469] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[470] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[471] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[472] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[473] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[474] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[475] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[476] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[477] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[478] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[479] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[480] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[481] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[482] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[483] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[484] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[485] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[486] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[487] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[488] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[489] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[490] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[491] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[492] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[493] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[494] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[495] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[496] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[497] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[498] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[499] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[500] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[501] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[502] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[503] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[504] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[505] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[506] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[507] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[508] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[509] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[510] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[511] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[512] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[513] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[514] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[515] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[516] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[517] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[518] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[519] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[520] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[521] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[522] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[523] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[524] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[525] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[526] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[527] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[528] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[529] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[530] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[531] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[532] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[533] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[534] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[535] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[536] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[537] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[538] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[539] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[540] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[541] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[542] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[543] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[544] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[545] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[546] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[547] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[548] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[549] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[550] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[551] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[552] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[553] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[554] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[555] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[556] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[557] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[558] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[559] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[560] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[561] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[562] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[563] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[564] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[565] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[566] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[567] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[568] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[569] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[570] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[571] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[572] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[573] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[574] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[575] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[576] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[577] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[578] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[579] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[580] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[581] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[582] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[583] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[584] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[585] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[586] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[587] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[588] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[589] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[590] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[591] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[592] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[593] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[594] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[595] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[596] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[597] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[598] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[599] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[600] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[601] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[602] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[603] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[604] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[605] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[606] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[607] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[608] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[609] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[610] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[611] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[612] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[613] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[614] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[615] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[616] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[617] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[618] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[619] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[620] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[621] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[622] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[623] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[624] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[625] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[626] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[627] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[628] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[629] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[630] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[631] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[632] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[633] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[634] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[635] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[636] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[637] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[638] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[639] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[640] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[641] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[642] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[643] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[644] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[645] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[646] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[647] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[648] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[649] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[650] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[651] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[652] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[653] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[654] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[655] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[656] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[657] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[658] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[659] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[660] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[661] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[662] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[663] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[664] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[665] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[666] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[667] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[668] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[669] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[670] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[671] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[672] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[673] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[674] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[675] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[676] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[677] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[678] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[679] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[680] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[681] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[682] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[683] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[684] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[685] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[686] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[687] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[688] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[689] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[690] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[691] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[692] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[693] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[694] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[695] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[696] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[697] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[698] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[699] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[700] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[701] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[702] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[703] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[704] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[705] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[706] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[707] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[708] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[709] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[710] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[711] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[712] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[713] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[714] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[715] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[716] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[717] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[718] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[719] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[720] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[721] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[722] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[723] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[724] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[725] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[726] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[727] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[728] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[729] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[730] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[731] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[732] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[733] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[734] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[735] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[736] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[737] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[738] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[739] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[740] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[741] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[742] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[743] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[744] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[745] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[746] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[747] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[748] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[749] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[750] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[751] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[752] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[753] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[754] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[755] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[756] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[757] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[758] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[759] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[760] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[761] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[762] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[763] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[764] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[765] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[766] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[767] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[768] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[769] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[770] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[771] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[772] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[773] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[774] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[775] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[776] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[777] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[778] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[779] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[780] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[781] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[782] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[783] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[784] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[785] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[786] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[787] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[788] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[789] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[790] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[791] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[792] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[793] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[794] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[795] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[796] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[797] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[798] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[799] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[800] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[801] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[802] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[803] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[804] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[805] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[806] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[807] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[808] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[809] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[810] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[811] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[812] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[813] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[814] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[815] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[816] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[817] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[818] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[819] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[820] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[821] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[822] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[823] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[824] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[825] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[826] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[827] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[828] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[829] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[830] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[831] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[832] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[833] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[834] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[835] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[836] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[837] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[838] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[839] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[840] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[841] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[842] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[843] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[844] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[845] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[846] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[847] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[848] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[849] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[850] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[851] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[852] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[853] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[854] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[855] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[856] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[857] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[858] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[859] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[860] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[861] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[862] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[863] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[864] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[865] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[866] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[867] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[868] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[869] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[870] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[871] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[872] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[873] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[874] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[875] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[876] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[877] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[878] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[879] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[880] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[881] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[882] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[883] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[884] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[885] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[886] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[887] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[888] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[889] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[890] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[891] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[892] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[893] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[894] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[895] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[896] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[897] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[898] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[899] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[900] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[901] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[902] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[903] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[904] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[905] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[906] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[907] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[908] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[909] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[910] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[911] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[912] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[913] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[914] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[915] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[916] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[917] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[918] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[919] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[920] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[921] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[922] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[923] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[924] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[925] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[926] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[927] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[928] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[929] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[930] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[931] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[932] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[933] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[934] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[935] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[936] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[937] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[938] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[939] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[940] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[941] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[942] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[943] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[944] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[945] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[946] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[947] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[948] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[949] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[950] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[951] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[952] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[953] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[954] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[955] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[956] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[957] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[958] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[959] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[960] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[961] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[962] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[963] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[964] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[965] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[966] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[967] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[968] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[969] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[970] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[971] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[972] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[973] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[974] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[975] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[976] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[977] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[978] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[979] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[980] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[981] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[982] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[983] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[984] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[985] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[986] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[987] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[988] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[989] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[990] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[991] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[992] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[993] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[994] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[995] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[996] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[997] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[998] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[999] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1000] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1001] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1002] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1003] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1004] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1005] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1006] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1007] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1008] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1009] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1010] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1011] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1012] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1013] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1014] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1015] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1016] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1017] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1018] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1019] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1020] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1021] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1022] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1023] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1024] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1025] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1026] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1027] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1028] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1029] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1030] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1031] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1032] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1033] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1034] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1035] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1036] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1037] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1038] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1039] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1040] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1041] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1042] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1043] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1044] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1045] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1046] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1047] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1048] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1049] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1050] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1051] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1052] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1053] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1054] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1055] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1056] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1057] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1058] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1059] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1060] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1061] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1062] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1063] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1064] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1065] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1066] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1067] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1068] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1069] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1070] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1071] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1072] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1073] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1074] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1075] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1076] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1077] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1078] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1079] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1080] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1081] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1082] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1083] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1084] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1085] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1086] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1087] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1088] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1089] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1090] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1091] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1092] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1093] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1094] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1095] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1096] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1097] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1098] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1099] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1100] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1101] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1102] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1103] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1104] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1105] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1106] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1107] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1108] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1109] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1110] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1111] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1112] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1113] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1114] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1115] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1116] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1117] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1118] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1119] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1120] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1121] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1122] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1123] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1124] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1125] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1126] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1127] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1128] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1129] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1130] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1131] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1132] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1133] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1134] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1135] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1136] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1137] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1138] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1139] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1140] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1141] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1142] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1143] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1144] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1145] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1146] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1147] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1148] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1149] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1150] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1151] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1152] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1153] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1154] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1155] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1156] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1157] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1158] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1159] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1160] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1161] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1162] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1163] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1164] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1165] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1166] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1167] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1168] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1169] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1170] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1171] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1172] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1173] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1174] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1175] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1176] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1177] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1178] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1179] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1180] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1181] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1182] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1183] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1184] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1185] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1186] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1187] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1188] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1189] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1190] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1191] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1192] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1193] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1194] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1195] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1196] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1197] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1198] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1199] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1200] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1201] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1202] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1203] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1204] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1205] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1206] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1207] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1208] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1209] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1210] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1211] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1212] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1213] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1214] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1215] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1216] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1217] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1218] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1219] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1220] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1221] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1222] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1223] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1224] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1225] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1226] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1227] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1228] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1229] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1230] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1231] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1232] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1233] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1234] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1235] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1236] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1237] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1238] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1239] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1240] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1241] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1242] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1243] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1244] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1245] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1246] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1247] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1248] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1249] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1250] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1251] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1252] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1253] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1254] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1255] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1256] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1257] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1258] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1259] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1260] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1261] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1262] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1263] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1264] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1265] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1266] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1267] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1268] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1269] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1270] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1271] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1272] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1273] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1274] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1275] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1276] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1277] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1278] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1279] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1280] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1281] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1282] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1283] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1284] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1285] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1286] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1287] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1288] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1289] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1290] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1291] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1292] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1293] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1294] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1295] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1296] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1297] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1298] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1299] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1300] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1301] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1302] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1303] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1304] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1305] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1306] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1307] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1308] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1309] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1310] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1311] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1312] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1313] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1314] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1315] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1316] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1317] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1318] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1319] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1320] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1321] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1322] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1323] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1324] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1325] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1326] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1327] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1328] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1329] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1330] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1331] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1332] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1333] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1334] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1335] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1336] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1337] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1338] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1339] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1340] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1341] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1342] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1343] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1344] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1345] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1346] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1347] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1348] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1349] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1350] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1351] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1352] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1353] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1354] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1355] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1356] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1357] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1358] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1359] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1360] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1361] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1362] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1363] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1364] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1365] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1366] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1367] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1368] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1369] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1370] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1371] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1372] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1373] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1374] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1375] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1376] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1377] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1378] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1379] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1380] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1381] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1382] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1383] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1384] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1385] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1386] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1387] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1388] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1389] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1390] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1391] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1392] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1393] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1394] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1395] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1396] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1397] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1398] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1399] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1400] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1401] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1402] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1403] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1404] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1405] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1406] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1407] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1408] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1409] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1410] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1411] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1412] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1413] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1414] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1415] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1416] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1417] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1418] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1419] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1420] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1421] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1422] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1423] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1424] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1425] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1426] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1427] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1428] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1429] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1430] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1431] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1432] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1433] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1434] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1435] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1436] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1437] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1438] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1439] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1440] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1441] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1442] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1443] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1444] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1445] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1446] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1447] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1448] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1449] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1450] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1451] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1452] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1453] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1454] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1455] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1456] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1457] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1458] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1459] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1460] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1461] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1462] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1463] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1464] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1465] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1466] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1467] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1468] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1469] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1470] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1471] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1472] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1473] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1474] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1475] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1476] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1477] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1478] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1479] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1480] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1481] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1482] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1483] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1484] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1485] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1486] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1487] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1488] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1489] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1490] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1491] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1492] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1493] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1494] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1495] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1496] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1497] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1498] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1499] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1500] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1501] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1502] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1503] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1504] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1505] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1506] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1507] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1508] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1509] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1510] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1511] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1512] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1513] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1514] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1515] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1516] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1517] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1518] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1519] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1520] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1521] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1522] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1523] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1524] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1525] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1526] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1527] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1528] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1529] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1530] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1531] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1532] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1533] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1534] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1535] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1536] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1537] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1538] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1539] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1540] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1541] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1542] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1543] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1544] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1545] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1546] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1547] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1548] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1549] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1550] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1551] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1552] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1553] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1554] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1555] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1556] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1557] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1558] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1559] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1560] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1561] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1562] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1563] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1564] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1565] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1566] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1567] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1568] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1569] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1570] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1571] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1572] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1573] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1574] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1575] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1576] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1577] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1578] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1579] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1580] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1581] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1582] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1583] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1584] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1585] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1586] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1587] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1588] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1589] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1590] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1591] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1592] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1593] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1594] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1595] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1596] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1597] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1598] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1599] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1600] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1601] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1602] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1603] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1604] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1605] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1606] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1607] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1608] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1609] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1610] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1611] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1612] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1613] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1614] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1615] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1616] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1617] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1618] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1619] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1620] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1621] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1622] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1623] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1624] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1625] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1626] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1627] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1628] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1629] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1630] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1631] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1632] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1633] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1634] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1635] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1636] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1637] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1638] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1639] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1640] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1641] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1642] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1643] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1644] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1645] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1646] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1647] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1648] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1649] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1650] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1651] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1652] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1653] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1654] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1655] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1656] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1657] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1658] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1659] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1660] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1661] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1662] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1663] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1664] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1665] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1666] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1667] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1668] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1669] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1670] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1671] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1672] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1673] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1674] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1675] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1676] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1677] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1678] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1679] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1680] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1681] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1682] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1683] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1684] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1685] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1686] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1687] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1688] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1689] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1690] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1691] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1692] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1693] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1694] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1695] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1696] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1697] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1698] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1699] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1700] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1701] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1702] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1703] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1704] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1705] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1706] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1707] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1708] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1709] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1710] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1711] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1712] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1713] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1714] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1715] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1716] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1717] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1718] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1719] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1720] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1721] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1722] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1723] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1724] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1725] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1726] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1727] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1728] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1729] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1730] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1731] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1732] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1733] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1734] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1735] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1736] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1737] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1738] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1739] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1740] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1741] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1742] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1743] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1744] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1745] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1746] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1747] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1748] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1749] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1750] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1751] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1752] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1753] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1754] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1755] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1756] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1757] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1758] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1759] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1760] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1761] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1762] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1763] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1764] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1765] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1766] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1767] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1768] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1769] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1770] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1771] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1772] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1773] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1774] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1775] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1776] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1777] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1778] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1779] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1780] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1781] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1782] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1783] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1784] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1785] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1786] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1787] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1788] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1789] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1790] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1791] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1792] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1793] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1794] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1795] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1796] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1797] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1798] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1799] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1800] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1801] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1802] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1803] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1804] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1805] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1806] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1807] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1808] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1809] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1810] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1811] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1812] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1813] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1814] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1815] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1816] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1817] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1818] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1819] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1820] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1821] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1822] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1823] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1824] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[1825] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[1826] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[1827] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[1828] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[1829] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[1830] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[1831] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[1832] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[1833] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[1834] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1835] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1836] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1837] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1838] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1839] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1840] = s[0] ? neg_SNs[24] : neg_SNs[24];
	assign level0[1841] = s[0] ? neg_SNs[24] : neg_SNs[24];
	assign level0[1842] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1843] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1844] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1845] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1846] = s[0] ? neg_SNs[28] : neg_SNs[28];
	assign level0[1847] = s[0] ? neg_SNs[28] : neg_SNs[28];
	assign level0[1848] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1849] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1850] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1851] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1852] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1853] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1854] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1855] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1856] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1857] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1858] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1859] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1860] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1861] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1862] = s[0] ? neg_SNs[37] : neg_SNs[37];
	assign level0[1863] = s[0] ? neg_SNs[37] : neg_SNs[37];
	assign level0[1864] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1865] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1866] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1867] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1868] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1869] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1870] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1871] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1872] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1873] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1874] = s[0] ? neg_SNs[56] : neg_SNs[56];
	assign level0[1875] = s[0] ? neg_SNs[56] : neg_SNs[56];
	assign level0[1876] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1877] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1878] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1879] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1880] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1881] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1882] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1883] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1884] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1885] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1886] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1887] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1888] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1889] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1890] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1891] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1892] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1893] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1894] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1895] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1896] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1897] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1898] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1899] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1900] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1901] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1902] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1903] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1904] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1905] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1906] = s[0] ? neg_SNs[92] : neg_SNs[92];
	assign level0[1907] = s[0] ? neg_SNs[92] : neg_SNs[92];
	assign level0[1908] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1909] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1910] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1911] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1912] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1913] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1914] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1915] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1916] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1917] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1918] = s[0] ? neg_SNs[111] : neg_SNs[111];
	assign level0[1919] = s[0] ? neg_SNs[111] : neg_SNs[111];
	assign level0[1920] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[1921] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[1922] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1923] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1924] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1925] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1926] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1927] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1928] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1929] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1930] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1931] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1932] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1933] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1934] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[1935] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[1936] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1937] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1938] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1939] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1940] = s[0] ? neg_SNs[124] : neg_SNs[124];
	assign level0[1941] = s[0] ? neg_SNs[124] : neg_SNs[124];
	assign level0[1942] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1943] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1944] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[1945] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[1946] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[1947] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[1948] = s[0] ? neg_SNs[132] : neg_SNs[132];
	assign level0[1949] = s[0] ? neg_SNs[132] : neg_SNs[132];
	assign level0[1950] = s[0] ? neg_SNs[14] : neg_SNs[14];
	assign level0[1951] = s[0] ? neg_SNs[15] : neg_SNs[15];
	assign level0[1952] = s[0] ? neg_SNs[17] : neg_SNs[17];
	assign level0[1953] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1954] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1955] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1956] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1957] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1958] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1959] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1960] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1961] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1962] = s[0] ? neg_SNs[40] : neg_SNs[40];
	assign level0[1963] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1964] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1965] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1966] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1967] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1968] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1969] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1970] = s[0] ? neg_SNs[54] : neg_SNs[54];
	assign level0[1971] = s[0] ? neg_SNs[56] : neg_SNs[56];
	assign level0[1972] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1973] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1974] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1975] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1976] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1977] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1978] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1979] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1980] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1981] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1982] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1983] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1984] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1985] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1986] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1987] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1988] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1989] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1990] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1991] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1992] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1993] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1994] = s[0] ? neg_SNs[92] : neg_SNs[92];
	assign level0[1995] = s[0] ? neg_SNs[94] : neg_SNs[94];
	assign level0[1996] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1997] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1998] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1999] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[2000] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[2001] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[2002] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[2003] = s[0] ? neg_SNs[108] : neg_SNs[108];
	assign level0[2004] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[2005] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[2006] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[2007] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[2008] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[2009] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[2010] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[2011] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2012] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2013] = s[0] ? neg_SNs[131] : neg_SNs[131];
	assign level0[2014] = s[0] ? neg_SNs[133] : neg_SNs[133];
	assign level0[2015] = s[0] ? neg_SNs[134] : neg_SNs[134];
	assign level0[2016] = s[0] ? pos_SNs[9] : pos_SNs[9];
	assign level0[2017] = s[0] ? pos_SNs[11] : pos_SNs[11];
	assign level0[2018] = s[0] ? neg_SNs[13] : neg_SNs[13];
	assign level0[2019] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[2020] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[2021] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[2022] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[2023] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[2024] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[2025] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[2026] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[2027] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[2028] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[2029] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[2030] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[2031] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[2032] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[2033] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[2034] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[2035] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[2036] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[2037] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[2038] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[2039] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[2040] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[2041] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[2042] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[2043] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[2044] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2045] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2046] = s[0] ? neg_SNs[135] : neg_SNs[135];
	assign level0[2047] = s[0] ? pos_SNs[138] : pos_SNs[138];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module hw_tree2  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[2] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[3] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[4] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[5] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[6] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[7] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[8] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[9] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[10] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[11] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[12] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[13] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[14] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[15] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[16] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[17] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[18] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[19] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[20] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[21] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[22] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[23] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[24] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[25] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[26] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[27] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[28] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[29] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[30] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[31] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[32] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[33] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[34] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[35] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[36] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[37] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[38] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[39] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[40] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[41] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[42] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[43] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[44] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[45] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[46] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[47] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[48] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[49] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[50] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[51] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[52] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[53] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[54] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[55] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[56] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[57] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[58] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[59] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[60] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[61] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[62] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[63] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[64] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[65] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[66] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[67] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[68] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[69] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[70] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[71] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[72] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[73] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[74] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[75] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[76] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[77] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[78] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[79] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[80] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[81] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[82] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[83] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[84] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[85] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[86] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[87] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[88] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[89] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[90] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[91] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[92] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[93] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[94] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[95] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[96] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[97] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[98] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[99] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[100] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[101] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[102] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[103] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[104] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[105] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[106] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[107] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[108] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[109] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[110] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[111] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[112] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[113] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[114] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[115] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[116] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[117] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[118] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[119] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[120] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[121] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[122] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[123] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[124] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[125] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[126] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[127] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[128] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[129] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[130] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[131] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[132] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[133] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[134] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[135] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[136] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[137] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[138] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[139] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[140] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[141] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[142] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[143] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[144] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[145] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[146] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[147] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[148] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[149] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[150] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[151] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[152] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[153] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[154] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[155] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[156] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[157] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[158] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[159] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[160] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[161] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[162] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[163] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[164] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[165] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[166] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[167] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[168] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[169] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[170] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[171] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[172] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[173] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[174] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[175] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[176] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[177] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[178] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[179] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[180] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[181] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[182] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[183] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[184] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[185] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[186] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[187] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[188] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[189] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[190] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[191] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[192] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[193] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[194] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[195] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[196] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[197] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[198] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[199] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[200] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[201] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[202] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[203] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[204] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[205] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[206] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[207] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[208] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[209] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[210] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[211] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[212] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[213] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[214] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[215] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[216] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[217] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[218] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[219] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[220] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[221] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[222] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[223] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[224] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[225] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[226] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[227] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[228] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[229] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[230] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[231] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[232] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[233] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[234] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[235] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[236] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[237] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[238] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[239] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[240] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[241] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[242] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[243] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[244] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[245] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[246] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[247] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[248] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[249] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[250] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[251] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[252] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[253] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[254] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[255] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[256] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[257] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[258] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[259] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[260] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[261] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[262] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[263] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[264] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[265] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[266] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[267] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[268] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[269] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[270] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[271] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[272] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[273] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[274] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[275] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[276] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[277] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[278] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[279] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[280] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[281] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[282] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[283] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[284] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[285] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[286] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[287] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[288] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[289] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[290] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[291] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[292] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[293] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[294] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[295] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[296] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[297] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[298] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[299] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[300] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[301] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[302] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[303] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[304] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[305] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[306] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[307] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[308] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[309] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[310] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[311] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[312] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[313] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[314] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[315] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[316] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[317] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[318] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[319] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[320] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[321] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[322] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[323] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[324] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[325] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[326] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[327] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[328] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[329] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[330] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[331] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[332] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[333] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[334] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[335] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[336] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[337] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[338] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[339] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[340] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[341] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[342] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[343] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[344] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[345] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[346] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[347] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[348] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[349] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[350] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[351] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[352] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[353] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[354] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[355] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[356] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[357] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[358] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[359] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[360] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[361] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[362] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[363] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[364] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[365] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[366] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[367] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[368] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[369] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[370] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[371] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[372] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[373] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[374] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[375] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[376] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[377] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[378] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[379] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[380] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[381] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[382] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[383] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[384] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[385] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[386] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[387] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[388] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[389] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[390] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[391] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[392] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[393] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[394] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[395] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[396] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[397] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[398] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[399] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[400] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[401] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[402] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[403] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[404] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[405] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[406] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[407] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[408] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[409] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[410] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[411] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[412] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[413] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[414] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[415] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[416] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[417] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[418] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[419] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[420] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[421] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[422] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[423] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[424] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[425] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[426] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[427] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[428] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[429] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[430] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[431] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[432] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[433] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[434] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[435] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[436] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[437] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[438] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[439] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[440] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[441] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[442] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[443] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[444] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[445] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[446] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[447] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[448] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[449] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[450] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[451] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[452] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[453] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[454] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[455] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[456] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[457] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[458] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[459] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[460] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[461] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[462] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[463] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[464] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[465] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[466] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[467] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[468] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[469] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[470] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[471] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[472] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[473] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[474] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[475] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[476] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[477] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[478] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[479] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[480] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[481] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[482] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[483] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[484] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[485] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[486] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[487] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[488] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[489] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[490] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[491] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[492] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[493] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[494] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[495] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[496] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[497] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[498] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[499] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[500] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[501] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[502] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[503] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[504] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[505] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[506] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[507] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[508] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[509] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[510] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[511] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[512] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[513] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[514] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[515] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[516] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[517] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[518] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[519] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[520] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[521] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[522] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[523] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[524] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[525] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[526] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[527] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[528] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[529] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[530] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[531] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[532] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[533] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[534] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[535] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[536] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[537] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[538] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[539] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[540] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[541] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[542] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[543] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[544] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[545] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[546] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[547] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[548] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[549] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[550] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[551] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[552] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[553] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[554] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[555] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[556] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[557] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[558] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[559] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[560] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[561] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[562] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[563] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[564] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[565] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[566] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[567] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[568] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[569] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[570] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[571] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[572] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[573] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[574] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[575] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[576] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[577] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[578] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[579] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[580] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[581] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[582] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[583] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[584] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[585] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[586] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[587] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[588] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[589] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[590] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[591] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[592] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[593] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[594] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[595] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[596] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[597] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[598] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[599] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[600] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[601] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[602] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[603] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[604] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[605] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[606] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[607] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[608] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[609] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[610] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[611] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[612] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[613] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[614] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[615] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[616] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[617] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[618] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[619] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[620] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[621] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[622] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[623] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[624] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[625] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[626] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[627] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[628] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[629] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[630] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[631] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[632] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[633] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[634] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[635] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[636] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[637] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[638] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[639] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[640] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[641] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[642] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[643] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[644] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[645] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[646] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[647] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[648] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[649] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[650] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[651] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[652] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[653] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[654] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[655] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[656] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[657] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[658] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[659] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[660] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[661] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[662] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[663] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[664] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[665] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[666] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[667] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[668] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[669] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[670] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[671] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[672] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[673] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[674] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[675] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[676] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[677] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[678] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[679] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[680] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[681] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[682] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[683] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[684] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[685] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[686] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[687] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[688] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[689] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[690] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[691] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[692] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[693] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[694] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[695] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[696] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[697] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[698] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[699] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[700] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[701] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[702] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[703] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[704] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[705] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[706] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[707] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[708] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[709] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[710] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[711] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[712] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[713] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[714] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[715] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[716] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[717] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[718] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[719] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[720] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[721] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[722] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[723] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[724] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[725] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[726] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[727] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[728] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[729] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[730] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[731] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[732] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[733] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[734] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[735] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[736] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[737] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[738] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[739] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[740] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[741] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[742] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[743] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[744] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[745] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[746] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[747] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[748] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[749] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[750] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[751] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[752] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[753] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[754] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[755] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[756] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[757] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[758] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[759] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[760] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[761] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[762] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[763] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[764] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[765] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[766] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[767] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[768] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[769] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[770] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[771] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[772] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[773] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[774] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[775] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[776] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[777] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[778] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[779] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[780] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[781] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[782] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[783] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[784] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[785] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[786] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[787] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[788] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[789] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[790] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[791] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[792] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[793] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[794] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[795] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[796] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[797] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[798] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[799] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[800] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[801] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[802] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[803] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[804] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[805] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[806] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[807] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[808] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[809] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[810] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[811] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[812] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[813] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[814] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[815] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[816] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[817] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[818] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[819] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[820] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[821] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[822] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[823] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[824] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[825] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[826] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[827] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[828] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[829] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[830] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[831] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[832] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[833] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[834] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[835] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[836] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[837] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[838] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[839] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[840] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[841] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[842] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[843] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[844] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[845] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[846] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[847] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[848] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[849] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[850] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[851] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[852] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[853] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[854] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[855] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[856] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[857] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[858] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[859] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[860] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[861] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[862] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[863] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[864] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[865] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[866] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[867] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[868] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[869] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[870] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[871] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[872] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[873] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[874] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[875] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[876] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[877] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[878] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[879] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[880] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[881] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[882] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[883] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[884] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[885] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[886] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[887] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[888] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[889] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[890] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[891] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[892] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[893] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[894] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[895] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[896] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[897] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[898] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[899] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[900] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[901] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[902] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[903] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[904] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[905] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[906] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[907] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[908] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[909] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[910] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[911] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[912] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[913] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[914] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[915] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[916] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[917] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[918] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[919] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[920] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[921] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[922] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[923] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[924] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[925] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[926] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[927] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[928] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[929] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[930] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[931] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[932] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[933] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[934] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[935] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[936] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[937] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[938] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[939] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[940] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[941] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[942] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[943] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[944] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[945] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[946] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[947] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[948] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[949] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[950] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[951] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[952] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[953] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[954] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[955] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[956] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[957] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[958] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[959] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[960] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[961] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[962] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[963] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[964] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[965] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[966] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[967] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[968] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[969] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[970] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[971] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[972] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[973] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[974] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[975] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[976] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[977] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[978] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[979] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[980] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[981] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[982] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[983] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[984] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[985] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[986] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[987] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[988] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[989] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[990] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[991] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[992] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[993] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[994] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[995] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[996] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[997] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[998] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[999] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1000] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1001] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1002] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1003] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1004] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1005] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1006] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1007] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1008] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1009] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1010] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1011] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1012] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1013] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1014] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1015] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1016] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1017] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1018] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1019] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1020] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1021] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1022] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1023] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1024] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1025] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1026] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1027] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1028] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1029] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1030] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1031] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1032] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1033] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1034] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1035] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1036] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1037] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1038] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1039] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1040] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1041] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1042] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1043] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1044] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1045] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1046] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1047] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1048] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1049] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1050] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1051] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1052] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1053] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1054] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1055] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1056] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1057] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1058] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1059] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1060] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1061] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1062] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1063] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1064] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1065] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1066] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1067] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1068] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1069] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1070] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1071] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1072] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1073] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1074] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1075] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1076] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1077] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1078] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1079] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1080] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1081] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1082] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1083] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1084] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1085] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1086] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1087] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1088] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1089] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1090] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1091] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1092] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1093] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1094] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1095] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1096] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1097] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1098] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1099] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1100] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1101] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1102] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1103] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1104] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1105] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1106] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1107] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1108] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1109] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1110] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1111] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1112] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1113] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1114] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1115] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1116] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1117] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1118] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1119] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1120] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1121] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1122] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1123] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1124] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1125] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1126] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1127] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1128] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1129] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1130] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1131] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1132] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1133] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1134] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1135] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1136] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1137] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1138] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1139] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1140] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1141] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1142] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1143] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1144] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1145] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1146] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1147] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1148] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1149] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1150] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1151] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1152] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1153] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1154] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1155] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1156] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1157] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1158] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1159] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1160] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1161] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1162] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1163] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1164] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1165] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1166] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1167] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1168] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1169] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1170] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1171] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1172] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1173] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1174] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1175] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1176] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1177] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1178] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1179] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1180] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1181] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1182] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1183] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1184] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1185] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1186] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1187] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1188] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1189] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1190] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1191] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1192] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1193] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1194] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1195] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1196] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1197] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1198] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1199] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1200] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1201] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1202] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1203] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1204] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1205] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1206] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1207] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1208] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1209] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1210] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1211] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1212] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1213] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1214] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1215] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1216] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1217] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1218] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1219] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1220] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1221] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1222] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1223] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1224] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1225] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1226] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1227] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1228] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1229] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1230] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1231] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1232] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1233] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1234] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1235] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1236] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1237] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1238] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1239] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1240] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1241] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1242] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1243] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1244] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1245] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1246] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1247] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1248] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1249] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1250] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1251] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1252] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1253] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1254] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1255] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1256] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1257] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1258] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1259] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1260] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1261] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1262] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1263] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1264] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1265] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1266] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1267] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1268] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1269] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1270] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1271] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1272] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1273] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1274] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1275] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1276] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1277] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1278] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1279] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1280] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1281] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1282] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1283] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1284] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1285] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1286] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1287] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1288] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1289] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1290] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1291] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1292] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1293] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1294] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1295] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1296] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1297] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1298] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1299] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1300] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1301] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1302] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1303] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1304] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1305] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1306] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1307] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1308] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1309] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1310] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1311] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1312] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1313] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1314] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1315] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1316] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1317] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1318] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1319] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1320] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1321] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1322] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1323] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1324] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1325] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1326] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1327] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1328] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1329] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1330] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1331] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1332] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1333] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1334] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1335] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1336] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1337] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1338] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1339] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1340] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1341] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1342] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1343] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1344] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1345] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1346] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1347] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1348] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1349] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1350] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1351] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1352] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1353] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1354] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1355] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1356] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1357] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1358] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1359] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1360] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1361] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1362] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1363] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1364] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1365] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1366] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1367] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1368] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1369] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1370] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1371] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1372] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1373] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1374] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1375] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1376] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1377] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1378] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1379] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1380] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1381] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1382] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1383] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1384] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1385] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1386] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1387] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1388] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1389] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1390] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1391] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1392] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1393] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1394] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1395] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1396] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1397] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1398] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1399] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1400] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1401] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1402] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1403] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1404] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1405] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1406] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1407] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1408] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1409] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1410] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1411] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1412] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1413] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1414] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1415] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1416] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1417] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1418] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1419] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1420] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1421] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1422] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1423] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1424] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1425] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1426] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1427] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1428] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1429] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1430] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1431] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1432] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1433] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1434] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1435] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1436] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1437] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1438] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1439] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1440] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1441] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1442] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1443] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1444] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1445] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1446] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1447] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1448] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1449] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1450] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1451] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1452] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1453] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1454] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1455] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1456] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1457] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1458] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1459] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1460] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1461] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1462] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1463] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1464] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1465] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1466] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1467] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1468] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1469] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1470] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1471] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1472] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1473] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1474] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1475] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1476] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1477] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1478] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1479] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1480] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1481] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1482] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1483] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1484] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1485] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1486] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1487] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1488] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1489] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1490] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1491] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1492] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1493] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1494] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1495] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1496] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1497] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1498] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1499] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1500] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1501] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1502] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1503] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1504] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1505] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1506] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1507] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1508] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1509] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1510] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1511] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1512] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1513] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1514] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1515] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1516] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1517] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1518] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1519] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1520] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1521] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1522] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1523] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1524] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1525] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1526] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1527] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1528] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1529] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1530] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1531] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1532] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1533] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1534] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1535] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1536] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1537] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1538] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1539] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1540] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1541] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1542] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1543] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1544] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1545] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1546] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1547] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1548] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1549] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1550] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1551] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1552] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1553] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1554] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1555] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1556] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1557] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1558] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1559] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1560] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1561] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1562] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1563] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1564] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1565] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1566] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1567] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1568] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1569] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1570] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1571] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1572] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1573] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1574] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1575] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1576] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1577] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1578] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1579] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1580] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1581] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1582] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1583] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1584] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1585] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1586] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1587] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1588] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1589] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1590] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1591] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1592] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1593] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1594] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1595] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1596] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1597] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1598] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1599] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1600] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1601] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1602] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1603] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1604] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1605] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1606] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1607] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1608] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1609] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1610] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1611] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1612] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1613] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1614] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1615] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1616] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1617] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1618] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1619] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1620] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1621] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1622] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1623] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1624] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1625] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1626] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1627] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1628] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1629] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1630] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1631] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1632] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1633] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1634] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1635] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1636] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1637] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1638] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1639] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1640] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1641] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1642] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1643] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1644] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1645] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1646] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1647] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1648] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1649] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1650] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1651] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1652] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1653] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1654] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1655] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1656] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1657] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1658] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1659] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1660] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1661] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1662] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1663] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1664] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1665] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1666] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1667] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1668] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1669] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1670] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1671] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1672] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[1673] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[1674] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[1675] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[1676] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1677] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1678] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1679] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1680] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1681] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1682] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1683] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1684] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1685] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1686] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1687] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1688] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1689] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1690] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1691] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1692] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1693] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1694] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1695] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1696] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1697] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1698] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1699] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1700] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1701] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1702] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1703] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1704] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1705] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1706] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1707] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1708] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1709] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1710] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1711] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1712] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1713] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1714] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1715] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1716] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1717] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1718] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1719] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1720] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1721] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1722] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1723] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1724] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1725] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1726] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1727] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1728] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1729] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1730] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1731] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1732] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1733] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1734] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1735] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1736] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1737] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1738] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1739] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1740] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1741] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1742] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1743] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1744] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1745] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1746] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1747] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1748] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1749] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1750] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1751] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1752] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1753] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1754] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1755] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1756] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1757] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1758] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1759] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1760] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1761] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1762] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1763] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1764] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1765] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1766] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1767] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1768] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1769] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1770] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1771] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1772] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1773] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1774] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1775] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1776] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1777] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1778] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1779] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1780] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1781] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1782] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1783] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1784] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1785] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1786] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1787] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1788] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1789] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1790] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1791] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1792] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1793] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1794] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1795] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1796] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1797] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1798] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1799] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1800] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1801] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1802] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1803] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1804] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1805] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1806] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1807] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1808] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1809] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1810] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1811] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1812] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1813] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1814] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1815] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1816] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1817] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1818] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1819] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1820] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1821] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1822] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1823] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1824] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1825] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1826] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1827] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1828] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1829] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1830] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1831] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1832] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1833] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1834] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1835] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1836] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1837] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1838] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1839] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1840] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1841] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1842] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1843] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[1844] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1845] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1846] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1847] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1848] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[1849] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[1850] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[1851] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[1852] = s[0] ? pos_SNs[16] : pos_SNs[16];
	assign level0[1853] = s[0] ? pos_SNs[16] : pos_SNs[16];
	assign level0[1854] = s[0] ? pos_SNs[17] : pos_SNs[17];
	assign level0[1855] = s[0] ? pos_SNs[17] : pos_SNs[17];
	assign level0[1856] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1857] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1858] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1859] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1860] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1861] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1862] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1863] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1864] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1865] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1866] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1867] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1868] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1869] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1870] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1871] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1872] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1873] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1874] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1875] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1876] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1877] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1878] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1879] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1880] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1881] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1882] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1883] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1884] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1885] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1886] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1887] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1888] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1889] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1890] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1891] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1892] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1893] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1894] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1895] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1896] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1897] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1898] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1899] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1900] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1901] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1902] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1903] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1904] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1905] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1906] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1907] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1908] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1909] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1910] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1911] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1912] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1913] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1914] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1915] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1916] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1917] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1918] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1919] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1920] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1921] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1922] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1923] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1924] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1925] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1926] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1927] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1928] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1929] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1930] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1931] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1932] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1933] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1934] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1935] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1936] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1937] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1938] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1939] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1940] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1941] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1942] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[1943] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[1944] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1945] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1946] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1947] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1948] = s[0] ? neg_SNs[128] : neg_SNs[128];
	assign level0[1949] = s[0] ? neg_SNs[128] : neg_SNs[128];
	assign level0[1950] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[1951] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[1952] = s[0] ? pos_SNs[131] : pos_SNs[131];
	assign level0[1953] = s[0] ? pos_SNs[131] : pos_SNs[131];
	assign level0[1954] = s[0] ? pos_SNs[132] : pos_SNs[132];
	assign level0[1955] = s[0] ? pos_SNs[132] : pos_SNs[132];
	assign level0[1956] = s[0] ? neg_SNs[13] : neg_SNs[13];
	assign level0[1957] = s[0] ? neg_SNs[14] : neg_SNs[14];
	assign level0[1958] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1959] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1960] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1961] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1962] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1963] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1964] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1965] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1966] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1967] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1968] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1969] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1970] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[1971] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1972] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1973] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1974] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1975] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1976] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1977] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1978] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1979] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1980] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1981] = s[0] ? neg_SNs[54] : neg_SNs[54];
	assign level0[1982] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[1983] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1984] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1985] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1986] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1987] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1988] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1989] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1990] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1991] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1992] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1993] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1994] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1995] = s[0] ? pos_SNs[93] : pos_SNs[93];
	assign level0[1996] = s[0] ? neg_SNs[94] : neg_SNs[94];
	assign level0[1997] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1998] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1999] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[2000] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[2001] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[2002] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[2003] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[2004] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[2005] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[2006] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[2007] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[2008] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[2009] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[2010] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[2011] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[2012] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[2013] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[2014] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[2015] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[2016] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[2017] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2018] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[2019] = s[0] ? neg_SNs[128] : neg_SNs[128];
	assign level0[2020] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[2021] = s[0] ? neg_SNs[134] : neg_SNs[134];
	assign level0[2022] = s[0] ? neg_SNs[135] : neg_SNs[135];
	assign level0[2023] = s[0] ? pos_SNs[10] : pos_SNs[10];
	assign level0[2024] = s[0] ? neg_SNs[12] : neg_SNs[12];
	assign level0[2025] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[2026] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[2027] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[2028] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[2029] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[2030] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[2031] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[2032] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[2033] = s[0] ? neg_SNs[54] : neg_SNs[54];
	assign level0[2034] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[2035] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[2036] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[2037] = s[0] ? neg_SNs[94] : neg_SNs[94];
	assign level0[2038] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[2039] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[2040] = s[0] ? pos_SNs[111] : pos_SNs[111];
	assign level0[2041] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[2042] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[2043] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[2044] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[2045] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2046] = s[0] ? pos_SNs[133] : pos_SNs[133];
	assign level0[2047] = s[0] ? pos_SNs[137] : pos_SNs[137];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module hw_tree3  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[2] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[3] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[4] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[5] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[6] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[7] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[8] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[9] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[10] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[11] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[12] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[13] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[14] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[15] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[16] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[17] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[18] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[19] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[20] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[21] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[22] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[23] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[24] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[25] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[26] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[27] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[28] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[29] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[30] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[31] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[32] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[33] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[34] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[35] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[36] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[37] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[38] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[39] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[40] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[41] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[42] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[43] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[44] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[45] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[46] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[47] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[48] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[49] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[50] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[51] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[52] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[53] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[54] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[55] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[56] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[57] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[58] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[59] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[60] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[61] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[62] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[63] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[64] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[65] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[66] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[67] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[68] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[69] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[70] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[71] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[72] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[73] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[74] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[75] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[76] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[77] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[78] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[79] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[80] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[81] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[82] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[83] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[84] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[85] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[86] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[87] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[88] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[89] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[90] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[91] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[92] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[93] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[94] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[95] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[96] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[97] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[98] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[99] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[100] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[101] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[102] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[103] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[104] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[105] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[106] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[107] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[108] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[109] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[110] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[111] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[112] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[113] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[114] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[115] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[116] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[117] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[118] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[119] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[120] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[121] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[122] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[123] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[124] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[125] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[126] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[127] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[128] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[129] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[130] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[131] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[132] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[133] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[134] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[135] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[136] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[137] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[138] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[139] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[140] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[141] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[142] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[143] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[144] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[145] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[146] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[147] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[148] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[149] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[150] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[151] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[152] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[153] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[154] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[155] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[156] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[157] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[158] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[159] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[160] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[161] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[162] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[163] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[164] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[165] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[166] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[167] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[168] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[169] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[170] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[171] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[172] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[173] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[174] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[175] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[176] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[177] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[178] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[179] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[180] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[181] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[182] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[183] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[184] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[185] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[186] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[187] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[188] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[189] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[190] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[191] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[192] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[193] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[194] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[195] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[196] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[197] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[198] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[199] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[200] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[201] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[202] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[203] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[204] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[205] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[206] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[207] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[208] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[209] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[210] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[211] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[212] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[213] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[214] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[215] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[216] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[217] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[218] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[219] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[220] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[221] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[222] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[223] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[224] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[225] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[226] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[227] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[228] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[229] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[230] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[231] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[232] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[233] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[234] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[235] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[236] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[237] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[238] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[239] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[240] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[241] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[242] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[243] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[244] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[245] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[246] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[247] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[248] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[249] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[250] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[251] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[252] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[253] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[254] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[255] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[256] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[257] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[258] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[259] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[260] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[261] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[262] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[263] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[264] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[265] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[266] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[267] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[268] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[269] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[270] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[271] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[272] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[273] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[274] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[275] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[276] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[277] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[278] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[279] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[280] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[281] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[282] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[283] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[284] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[285] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[286] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[287] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[288] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[289] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[290] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[291] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[292] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[293] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[294] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[295] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[296] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[297] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[298] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[299] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[300] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[301] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[302] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[303] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[304] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[305] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[306] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[307] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[308] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[309] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[310] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[311] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[312] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[313] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[314] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[315] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[316] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[317] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[318] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[319] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[320] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[321] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[322] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[323] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[324] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[325] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[326] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[327] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[328] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[329] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[330] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[331] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[332] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[333] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[334] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[335] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[336] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[337] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[338] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[339] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[340] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[341] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[342] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[343] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[344] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[345] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[346] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[347] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[348] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[349] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[350] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[351] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[352] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[353] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[354] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[355] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[356] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[357] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[358] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[359] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[360] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[361] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[362] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[363] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[364] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[365] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[366] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[367] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[368] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[369] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[370] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[371] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[372] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[373] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[374] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[375] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[376] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[377] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[378] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[379] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[380] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[381] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[382] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[383] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[384] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[385] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[386] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[387] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[388] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[389] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[390] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[391] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[392] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[393] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[394] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[395] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[396] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[397] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[398] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[399] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[400] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[401] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[402] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[403] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[404] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[405] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[406] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[407] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[408] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[409] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[410] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[411] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[412] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[413] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[414] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[415] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[416] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[417] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[418] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[419] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[420] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[421] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[422] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[423] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[424] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[425] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[426] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[427] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[428] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[429] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[430] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[431] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[432] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[433] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[434] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[435] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[436] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[437] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[438] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[439] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[440] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[441] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[442] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[443] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[444] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[445] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[446] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[447] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[448] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[449] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[450] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[451] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[452] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[453] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[454] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[455] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[456] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[457] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[458] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[459] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[460] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[461] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[462] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[463] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[464] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[465] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[466] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[467] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[468] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[469] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[470] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[471] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[472] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[473] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[474] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[475] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[476] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[477] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[478] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[479] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[480] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[481] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[482] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[483] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[484] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[485] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[486] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[487] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[488] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[489] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[490] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[491] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[492] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[493] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[494] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[495] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[496] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[497] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[498] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[499] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[500] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[501] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[502] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[503] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[504] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[505] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[506] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[507] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[508] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[509] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[510] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[511] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[512] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[513] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[514] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[515] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[516] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[517] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[518] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[519] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[520] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[521] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[522] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[523] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[524] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[525] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[526] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[527] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[528] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[529] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[530] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[531] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[532] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[533] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[534] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[535] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[536] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[537] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[538] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[539] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[540] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[541] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[542] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[543] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[544] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[545] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[546] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[547] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[548] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[549] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[550] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[551] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[552] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[553] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[554] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[555] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[556] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[557] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[558] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[559] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[560] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[561] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[562] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[563] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[564] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[565] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[566] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[567] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[568] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[569] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[570] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[571] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[572] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[573] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[574] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[575] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[576] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[577] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[578] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[579] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[580] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[581] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[582] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[583] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[584] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[585] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[586] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[587] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[588] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[589] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[590] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[591] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[592] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[593] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[594] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[595] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[596] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[597] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[598] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[599] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[600] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[601] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[602] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[603] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[604] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[605] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[606] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[607] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[608] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[609] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[610] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[611] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[612] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[613] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[614] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[615] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[616] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[617] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[618] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[619] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[620] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[621] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[622] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[623] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[624] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[625] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[626] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[627] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[628] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[629] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[630] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[631] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[632] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[633] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[634] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[635] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[636] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[637] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[638] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[639] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[640] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[641] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[642] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[643] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[644] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[645] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[646] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[647] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[648] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[649] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[650] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[651] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[652] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[653] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[654] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[655] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[656] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[657] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[658] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[659] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[660] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[661] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[662] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[663] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[664] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[665] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[666] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[667] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[668] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[669] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[670] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[671] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[672] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[673] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[674] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[675] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[676] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[677] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[678] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[679] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[680] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[681] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[682] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[683] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[684] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[685] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[686] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[687] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[688] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[689] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[690] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[691] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[692] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[693] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[694] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[695] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[696] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[697] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[698] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[699] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[700] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[701] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[702] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[703] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[704] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[705] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[706] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[707] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[708] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[709] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[710] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[711] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[712] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[713] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[714] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[715] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[716] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[717] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[718] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[719] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[720] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[721] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[722] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[723] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[724] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[725] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[726] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[727] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[728] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[729] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[730] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[731] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[732] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[733] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[734] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[735] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[736] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[737] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[738] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[739] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[740] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[741] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[742] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[743] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[744] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[745] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[746] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[747] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[748] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[749] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[750] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[751] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[752] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[753] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[754] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[755] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[756] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[757] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[758] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[759] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[760] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[761] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[762] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[763] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[764] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[765] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[766] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[767] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[768] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[769] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[770] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[771] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[772] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[773] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[774] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[775] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[776] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[777] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[778] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[779] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[780] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[781] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[782] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[783] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[784] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[785] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[786] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[787] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[788] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[789] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[790] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[791] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[792] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[793] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[794] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[795] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[796] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[797] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[798] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[799] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[800] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[801] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[802] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[803] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[804] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[805] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[806] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[807] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[808] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[809] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[810] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[811] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[812] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[813] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[814] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[815] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[816] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[817] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[818] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[819] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[820] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[821] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[822] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[823] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[824] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[825] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[826] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[827] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[828] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[829] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[830] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[831] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[832] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[833] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[834] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[835] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[836] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[837] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[838] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[839] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[840] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[841] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[842] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[843] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[844] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[845] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[846] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[847] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[848] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[849] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[850] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[851] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[852] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[853] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[854] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[855] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[856] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[857] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[858] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[859] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[860] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[861] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[862] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[863] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[864] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[865] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[866] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[867] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[868] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[869] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[870] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[871] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[872] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[873] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[874] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[875] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[876] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[877] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[878] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[879] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[880] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[881] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[882] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[883] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[884] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[885] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[886] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[887] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[888] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[889] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[890] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[891] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[892] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[893] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[894] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[895] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[896] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[897] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[898] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[899] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[900] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[901] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[902] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[903] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[904] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[905] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[906] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[907] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[908] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[909] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[910] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[911] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[912] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[913] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[914] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[915] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[916] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[917] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[918] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[919] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[920] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[921] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[922] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[923] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[924] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[925] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[926] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[927] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[928] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[929] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[930] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[931] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[932] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[933] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[934] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[935] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[936] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[937] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[938] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[939] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[940] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[941] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[942] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[943] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[944] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[945] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[946] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[947] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[948] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[949] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[950] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[951] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[952] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[953] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[954] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[955] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[956] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[957] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[958] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[959] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[960] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[961] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[962] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[963] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[964] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[965] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[966] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[967] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[968] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[969] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[970] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[971] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[972] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[973] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[974] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[975] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[976] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[977] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[978] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[979] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[980] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[981] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[982] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[983] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[984] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[985] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[986] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[987] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[988] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[989] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[990] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[991] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[992] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[993] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[994] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[995] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[996] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[997] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[998] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[999] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1000] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1001] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1002] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1003] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1004] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1005] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1006] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1007] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1008] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1009] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1010] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1011] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1012] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1013] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1014] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1015] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1016] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1017] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1018] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1019] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1020] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1021] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1022] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1023] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1024] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1025] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1026] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1027] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1028] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1029] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1030] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1031] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1032] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1033] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1034] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1035] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1036] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1037] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1038] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1039] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1040] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1041] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1042] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1043] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1044] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1045] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1046] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1047] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1048] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1049] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1050] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1051] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1052] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1053] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1054] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1055] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1056] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1057] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1058] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1059] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1060] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1061] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1062] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1063] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1064] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1065] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1066] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1067] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1068] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1069] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1070] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1071] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1072] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1073] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1074] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1075] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1076] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1077] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1078] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1079] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1080] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1081] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1082] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1083] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1084] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1085] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1086] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1087] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1088] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1089] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1090] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1091] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1092] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1093] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1094] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1095] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1096] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1097] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1098] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1099] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1100] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1101] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1102] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1103] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1104] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1105] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1106] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1107] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1108] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1109] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1110] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1111] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1112] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1113] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1114] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1115] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1116] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1117] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1118] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1119] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1120] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1121] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1122] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1123] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1124] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1125] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1126] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1127] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1128] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1129] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1130] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1131] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1132] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1133] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1134] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1135] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1136] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1137] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1138] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1139] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1140] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1141] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1142] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1143] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1144] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1145] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1146] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1147] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1148] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1149] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1150] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1151] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1152] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1153] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1154] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1155] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1156] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1157] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1158] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1159] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1160] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1161] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1162] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1163] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1164] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1165] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1166] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1167] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1168] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1169] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1170] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1171] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1172] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1173] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1174] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1175] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1176] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1177] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1178] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1179] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1180] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1181] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1182] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1183] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1184] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1185] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1186] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1187] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1188] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1189] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1190] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1191] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1192] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1193] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1194] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1195] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1196] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1197] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1198] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1199] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1200] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1201] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1202] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1203] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1204] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1205] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1206] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1207] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1208] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1209] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1210] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1211] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1212] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1213] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1214] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1215] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1216] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1217] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1218] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1219] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1220] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1221] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1222] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1223] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1224] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1225] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1226] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1227] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1228] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1229] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1230] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1231] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1232] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1233] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1234] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1235] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1236] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1237] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1238] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1239] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1240] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1241] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1242] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1243] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1244] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1245] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1246] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1247] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1248] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1249] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1250] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1251] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1252] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1253] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1254] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1255] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1256] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1257] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1258] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1259] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1260] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1261] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1262] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1263] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1264] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1265] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1266] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1267] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1268] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1269] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1270] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1271] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1272] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1273] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1274] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1275] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1276] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1277] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1278] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1279] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1280] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1281] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1282] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1283] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1284] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1285] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1286] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1287] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1288] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1289] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1290] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1291] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1292] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1293] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1294] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1295] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1296] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1297] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1298] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1299] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1300] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1301] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1302] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1303] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1304] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1305] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1306] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1307] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1308] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1309] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1310] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1311] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1312] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1313] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1314] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1315] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1316] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1317] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1318] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1319] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1320] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1321] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1322] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1323] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1324] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1325] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1326] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1327] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1328] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1329] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1330] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1331] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1332] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1333] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1334] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1335] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1336] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1337] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1338] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1339] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1340] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1341] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1342] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1343] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1344] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1345] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1346] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1347] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1348] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1349] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1350] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1351] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1352] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1353] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1354] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1355] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1356] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1357] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1358] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1359] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1360] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1361] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1362] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1363] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1364] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1365] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1366] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1367] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1368] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1369] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1370] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1371] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1372] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1373] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1374] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1375] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1376] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1377] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1378] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1379] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1380] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1381] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1382] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1383] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1384] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1385] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1386] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1387] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1388] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1389] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1390] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1391] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1392] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1393] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1394] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1395] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1396] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1397] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1398] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1399] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1400] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1401] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1402] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1403] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1404] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1405] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1406] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1407] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1408] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1409] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1410] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1411] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1412] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1413] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1414] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1415] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1416] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1417] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1418] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1419] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1420] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1421] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1422] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1423] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1424] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1425] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1426] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1427] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1428] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1429] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1430] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1431] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1432] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1433] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1434] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1435] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1436] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1437] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1438] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1439] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1440] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1441] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1442] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1443] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1444] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1445] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1446] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1447] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1448] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1449] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1450] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1451] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1452] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1453] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1454] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1455] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1456] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1457] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1458] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1459] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1460] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1461] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1462] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1463] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1464] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1465] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1466] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1467] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1468] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1469] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1470] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1471] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1472] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1473] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1474] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1475] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1476] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1477] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1478] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1479] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1480] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1481] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1482] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1483] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1484] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1485] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1486] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1487] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1488] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1489] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1490] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1491] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1492] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1493] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1494] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1495] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1496] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1497] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1498] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1499] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1500] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1501] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1502] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1503] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1504] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1505] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1506] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1507] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1508] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1509] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1510] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1511] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1512] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1513] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1514] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1515] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1516] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1517] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1518] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1519] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1520] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1521] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1522] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1523] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1524] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1525] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1526] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1527] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1528] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1529] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1530] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1531] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1532] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1533] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1534] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1535] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1536] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1537] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1538] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1539] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1540] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1541] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1542] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1543] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1544] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1545] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1546] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1547] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1548] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1549] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1550] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1551] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1552] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1553] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1554] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1555] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1556] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1557] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1558] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1559] = s[0] ? pos_SNs[73] : pos_SNs[73];
	assign level0[1560] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1561] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1562] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1563] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1564] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1565] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1566] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1567] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1568] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1569] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1570] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1571] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1572] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1573] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1574] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1575] = s[0] ? pos_SNs[75] : pos_SNs[75];
	assign level0[1576] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1577] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1578] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1579] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1580] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1581] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1582] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1583] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1584] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1585] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1586] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1587] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1588] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1589] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1590] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1591] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1592] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1593] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1594] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1595] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1596] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1597] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1598] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1599] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1600] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1601] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1602] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1603] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1604] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1605] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1606] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1607] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1608] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1609] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1610] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1611] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1612] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1613] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1614] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1615] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1616] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1617] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1618] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1619] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1620] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1621] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1622] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1623] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1624] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1625] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1626] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1627] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1628] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1629] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1630] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1631] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1632] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1633] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1634] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1635] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1636] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1637] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1638] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1639] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1640] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1641] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1642] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1643] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1644] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1645] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1646] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1647] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1648] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1649] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1650] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1651] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1652] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1653] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1654] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1655] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1656] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1657] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1658] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1659] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1660] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1661] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1662] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1663] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1664] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1665] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1666] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1667] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1668] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1669] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1670] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1671] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1672] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1673] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1674] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1675] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1676] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1677] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1678] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1679] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1680] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1681] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1682] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1683] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1684] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1685] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1686] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1687] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1688] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1689] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1690] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1691] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1692] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1693] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1694] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1695] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1696] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1697] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1698] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1699] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1700] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1701] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1702] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1703] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1704] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1705] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1706] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1707] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1708] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1709] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1710] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1711] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1712] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1713] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1714] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1715] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1716] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1717] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1718] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1719] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1720] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1721] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1722] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1723] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1724] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1725] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1726] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1727] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1728] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1729] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1730] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1731] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1732] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1733] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1734] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1735] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1736] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1737] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1738] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1739] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1740] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1741] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1742] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1743] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1744] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1745] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1746] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1747] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1748] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1749] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1750] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1751] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1752] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1753] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1754] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1755] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1756] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1757] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1758] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1759] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1760] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1761] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1762] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1763] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1764] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1765] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1766] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1767] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1768] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1769] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1770] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1771] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1772] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1773] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1774] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1775] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1776] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1777] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1778] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1779] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1780] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1781] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1782] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1783] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1784] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1785] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1786] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1787] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1788] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1789] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1790] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1791] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1792] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1793] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1794] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1795] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1796] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1797] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1798] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1799] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1800] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1801] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1802] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1803] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1804] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1805] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1806] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1807] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1808] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1809] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1810] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1811] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1812] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1813] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1814] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1815] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1816] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1817] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1818] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1819] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1820] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1821] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1822] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1823] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1824] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1825] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1826] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1827] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1828] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1829] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1830] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1831] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1832] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1833] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1834] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1835] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1836] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1837] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1838] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1839] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1840] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1841] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1842] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1843] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1844] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1845] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1846] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1847] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1848] = s[0] ? neg_SNs[17] : neg_SNs[17];
	assign level0[1849] = s[0] ? neg_SNs[17] : neg_SNs[17];
	assign level0[1850] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1851] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1852] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1853] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1854] = s[0] ? neg_SNs[22] : neg_SNs[22];
	assign level0[1855] = s[0] ? neg_SNs[22] : neg_SNs[22];
	assign level0[1856] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1857] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1858] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1859] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1860] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1861] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1862] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1863] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1864] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1865] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1866] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1867] = s[0] ? neg_SNs[43] : neg_SNs[43];
	assign level0[1868] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1869] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1870] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1871] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1872] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1873] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1874] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1875] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1876] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1877] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1878] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1879] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1880] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1881] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1882] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1883] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1884] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1885] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1886] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1887] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1888] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1889] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1890] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1891] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1892] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1893] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1894] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1895] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1896] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1897] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1898] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1899] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1900] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1901] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1902] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1903] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1904] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1905] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1906] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1907] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1908] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1909] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1910] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1911] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1912] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1913] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1914] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1915] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1916] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1917] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1918] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1919] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1920] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1921] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1922] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1923] = s[0] ? neg_SNs[105] : neg_SNs[105];
	assign level0[1924] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1925] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1926] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1927] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1928] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1929] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1930] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1931] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1932] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[1933] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[1934] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[1935] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[1936] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[1937] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[1938] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[1939] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[1940] = s[0] ? neg_SNs[131] : neg_SNs[131];
	assign level0[1941] = s[0] ? neg_SNs[131] : neg_SNs[131];
	assign level0[1942] = s[0] ? pos_SNs[14] : pos_SNs[14];
	assign level0[1943] = s[0] ? pos_SNs[15] : pos_SNs[15];
	assign level0[1944] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[1945] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1946] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1947] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1948] = s[0] ? neg_SNs[22] : neg_SNs[22];
	assign level0[1949] = s[0] ? pos_SNs[23] : pos_SNs[23];
	assign level0[1950] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1951] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[1952] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[1953] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1954] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1955] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1956] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1957] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1958] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[1959] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1960] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1961] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1962] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1963] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1964] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1965] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1966] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1967] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1968] = s[0] ? neg_SNs[59] : neg_SNs[59];
	assign level0[1969] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1970] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1971] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1972] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1973] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1974] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1975] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1976] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1977] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1978] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1979] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1980] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1981] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1982] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1983] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1984] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1985] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1986] = s[0] ? neg_SNs[89] : neg_SNs[89];
	assign level0[1987] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1988] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1989] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1990] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1991] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1992] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1993] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1994] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1995] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1996] = s[0] ? pos_SNs[109] : pos_SNs[109];
	assign level0[1997] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[1998] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1999] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[2000] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[2001] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[2002] = s[0] ? neg_SNs[121] : neg_SNs[121];
	assign level0[2003] = s[0] ? neg_SNs[123] : neg_SNs[123];
	assign level0[2004] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[2005] = s[0] ? pos_SNs[125] : pos_SNs[125];
	assign level0[2006] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[2007] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[2008] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2009] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[2010] = s[0] ? neg_SNs[132] : neg_SNs[132];
	assign level0[2011] = s[0] ? pos_SNs[133] : pos_SNs[133];
	assign level0[2012] = s[0] ? pos_SNs[134] : pos_SNs[134];
	assign level0[2013] = s[0] ? pos_SNs[10] : pos_SNs[10];
	assign level0[2014] = s[0] ? neg_SNs[13] : neg_SNs[13];
	assign level0[2015] = s[0] ? neg_SNs[17] : neg_SNs[17];
	assign level0[2016] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[2017] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[2018] = s[0] ? neg_SNs[27] : neg_SNs[27];
	assign level0[2019] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[2020] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[2021] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[2022] = s[0] ? pos_SNs[39] : pos_SNs[39];
	assign level0[2023] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[2024] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[2025] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[2026] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[2027] = s[0] ? pos_SNs[55] : pos_SNs[55];
	assign level0[2028] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[2029] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[2030] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[2031] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[2032] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[2033] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[2034] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[2035] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[2036] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[2037] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[2038] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[2039] = s[0] ? neg_SNs[110] : neg_SNs[110];
	assign level0[2040] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[2041] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[2042] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[2043] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[2044] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[2045] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2046] = s[0] ? pos_SNs[133] : pos_SNs[133];
	assign level0[2047] = s[0] ? neg_SNs[136] : neg_SNs[136];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module hw_tree4  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[2] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[3] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[4] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[5] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[6] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[7] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[8] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[9] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[10] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[11] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[12] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[13] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[14] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[15] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[16] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[17] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[18] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[19] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[20] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[21] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[22] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[23] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[24] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[25] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[26] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[27] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[28] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[29] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[30] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[31] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[32] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[33] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[34] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[35] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[36] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[37] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[38] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[39] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[40] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[41] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[42] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[43] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[44] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[45] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[46] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[47] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[48] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[49] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[50] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[51] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[52] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[53] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[54] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[55] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[56] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[57] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[58] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[59] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[60] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[61] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[62] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[63] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[64] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[65] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[66] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[67] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[68] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[69] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[70] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[71] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[72] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[73] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[74] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[75] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[76] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[77] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[78] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[79] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[80] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[81] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[82] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[83] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[84] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[85] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[86] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[87] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[88] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[89] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[90] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[91] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[92] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[93] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[94] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[95] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[96] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[97] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[98] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[99] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[100] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[101] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[102] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[103] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[104] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[105] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[106] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[107] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[108] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[109] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[110] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[111] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[112] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[113] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[114] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[115] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[116] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[117] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[118] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[119] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[120] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[121] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[122] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[123] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[124] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[125] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[126] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[127] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[128] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[129] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[130] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[131] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[132] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[133] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[134] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[135] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[136] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[137] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[138] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[139] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[140] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[141] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[142] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[143] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[144] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[145] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[146] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[147] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[148] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[149] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[150] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[151] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[152] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[153] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[154] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[155] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[156] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[157] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[158] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[159] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[160] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[161] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[162] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[163] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[164] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[165] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[166] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[167] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[168] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[169] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[170] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[171] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[172] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[173] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[174] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[175] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[176] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[177] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[178] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[179] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[180] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[181] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[182] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[183] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[184] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[185] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[186] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[187] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[188] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[189] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[190] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[191] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[192] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[193] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[194] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[195] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[196] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[197] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[198] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[199] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[200] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[201] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[202] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[203] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[204] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[205] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[206] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[207] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[208] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[209] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[210] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[211] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[212] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[213] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[214] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[215] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[216] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[217] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[218] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[219] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[220] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[221] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[222] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[223] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[224] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[225] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[226] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[227] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[228] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[229] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[230] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[231] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[232] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[233] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[234] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[235] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[236] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[237] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[238] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[239] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[240] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[241] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[242] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[243] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[244] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[245] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[246] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[247] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[248] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[249] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[250] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[251] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[252] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[253] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[254] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[255] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[256] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[257] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[258] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[259] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[260] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[261] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[262] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[263] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[264] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[265] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[266] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[267] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[268] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[269] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[270] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[271] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[272] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[273] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[274] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[275] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[276] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[277] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[278] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[279] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[280] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[281] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[282] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[283] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[284] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[285] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[286] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[287] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[288] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[289] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[290] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[291] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[292] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[293] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[294] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[295] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[296] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[297] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[298] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[299] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[300] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[301] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[302] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[303] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[304] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[305] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[306] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[307] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[308] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[309] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[310] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[311] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[312] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[313] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[314] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[315] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[316] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[317] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[318] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[319] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[320] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[321] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[322] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[323] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[324] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[325] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[326] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[327] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[328] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[329] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[330] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[331] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[332] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[333] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[334] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[335] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[336] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[337] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[338] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[339] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[340] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[341] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[342] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[343] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[344] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[345] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[346] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[347] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[348] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[349] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[350] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[351] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[352] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[353] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[354] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[355] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[356] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[357] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[358] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[359] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[360] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[361] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[362] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[363] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[364] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[365] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[366] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[367] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[368] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[369] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[370] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[371] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[372] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[373] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[374] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[375] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[376] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[377] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[378] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[379] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[380] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[381] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[382] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[383] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[384] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[385] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[386] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[387] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[388] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[389] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[390] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[391] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[392] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[393] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[394] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[395] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[396] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[397] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[398] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[399] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[400] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[401] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[402] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[403] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[404] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[405] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[406] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[407] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[408] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[409] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[410] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[411] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[412] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[413] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[414] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[415] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[416] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[417] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[418] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[419] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[420] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[421] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[422] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[423] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[424] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[425] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[426] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[427] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[428] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[429] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[430] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[431] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[432] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[433] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[434] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[435] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[436] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[437] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[438] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[439] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[440] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[441] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[442] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[443] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[444] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[445] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[446] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[447] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[448] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[449] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[450] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[451] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[452] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[453] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[454] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[455] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[456] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[457] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[458] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[459] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[460] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[461] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[462] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[463] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[464] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[465] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[466] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[467] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[468] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[469] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[470] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[471] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[472] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[473] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[474] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[475] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[476] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[477] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[478] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[479] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[480] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[481] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[482] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[483] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[484] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[485] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[486] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[487] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[488] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[489] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[490] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[491] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[492] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[493] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[494] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[495] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[496] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[497] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[498] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[499] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[500] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[501] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[502] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[503] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[504] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[505] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[506] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[507] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[508] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[509] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[510] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[511] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[512] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[513] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[514] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[515] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[516] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[517] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[518] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[519] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[520] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[521] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[522] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[523] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[524] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[525] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[526] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[527] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[528] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[529] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[530] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[531] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[532] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[533] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[534] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[535] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[536] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[537] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[538] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[539] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[540] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[541] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[542] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[543] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[544] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[545] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[546] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[547] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[548] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[549] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[550] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[551] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[552] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[553] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[554] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[555] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[556] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[557] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[558] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[559] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[560] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[561] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[562] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[563] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[564] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[565] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[566] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[567] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[568] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[569] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[570] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[571] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[572] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[573] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[574] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[575] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[576] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[577] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[578] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[579] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[580] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[581] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[582] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[583] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[584] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[585] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[586] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[587] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[588] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[589] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[590] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[591] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[592] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[593] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[594] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[595] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[596] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[597] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[598] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[599] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[600] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[601] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[602] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[603] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[604] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[605] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[606] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[607] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[608] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[609] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[610] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[611] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[612] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[613] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[614] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[615] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[616] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[617] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[618] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[619] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[620] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[621] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[622] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[623] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[624] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[625] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[626] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[627] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[628] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[629] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[630] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[631] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[632] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[633] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[634] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[635] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[636] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[637] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[638] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[639] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[640] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[641] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[642] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[643] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[644] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[645] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[646] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[647] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[648] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[649] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[650] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[651] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[652] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[653] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[654] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[655] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[656] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[657] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[658] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[659] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[660] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[661] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[662] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[663] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[664] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[665] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[666] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[667] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[668] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[669] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[670] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[671] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[672] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[673] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[674] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[675] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[676] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[677] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[678] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[679] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[680] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[681] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[682] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[683] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[684] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[685] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[686] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[687] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[688] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[689] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[690] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[691] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[692] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[693] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[694] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[695] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[696] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[697] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[698] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[699] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[700] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[701] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[702] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[703] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[704] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[705] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[706] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[707] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[708] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[709] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[710] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[711] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[712] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[713] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[714] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[715] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[716] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[717] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[718] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[719] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[720] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[721] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[722] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[723] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[724] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[725] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[726] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[727] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[728] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[729] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[730] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[731] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[732] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[733] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[734] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[735] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[736] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[737] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[738] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[739] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[740] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[741] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[742] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[743] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[744] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[745] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[746] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[747] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[748] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[749] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[750] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[751] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[752] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[753] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[754] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[755] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[756] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[757] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[758] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[759] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[760] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[761] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[762] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[763] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[764] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[765] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[766] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[767] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[768] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[769] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[770] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[771] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[772] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[773] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[774] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[775] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[776] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[777] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[778] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[779] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[780] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[781] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[782] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[783] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[784] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[785] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[786] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[787] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[788] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[789] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[790] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[791] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[792] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[793] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[794] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[795] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[796] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[797] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[798] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[799] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[800] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[801] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[802] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[803] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[804] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[805] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[806] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[807] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[808] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[809] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[810] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[811] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[812] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[813] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[814] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[815] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[816] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[817] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[818] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[819] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[820] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[821] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[822] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[823] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[824] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[825] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[826] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[827] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[828] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[829] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[830] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[831] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[832] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[833] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[834] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[835] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[836] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[837] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[838] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[839] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[840] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[841] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[842] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[843] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[844] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[845] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[846] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[847] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[848] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[849] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[850] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[851] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[852] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[853] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[854] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[855] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[856] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[857] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[858] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[859] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[860] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[861] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[862] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[863] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[864] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[865] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[866] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[867] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[868] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[869] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[870] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[871] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[872] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[873] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[874] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[875] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[876] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[877] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[878] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[879] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[880] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[881] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[882] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[883] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[884] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[885] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[886] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[887] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[888] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[889] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[890] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[891] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[892] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[893] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[894] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[895] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[896] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[897] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[898] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[899] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[900] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[901] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[902] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[903] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[904] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[905] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[906] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[907] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[908] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[909] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[910] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[911] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[912] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[913] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[914] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[915] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[916] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[917] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[918] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[919] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[920] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[921] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[922] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[923] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[924] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[925] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[926] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[927] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[928] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[929] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[930] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[931] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[932] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[933] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[934] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[935] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[936] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[937] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[938] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[939] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[940] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[941] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[942] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[943] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[944] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[945] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[946] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[947] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[948] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[949] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[950] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[951] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[952] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[953] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[954] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[955] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[956] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[957] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[958] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[959] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[960] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[961] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[962] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[963] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[964] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[965] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[966] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[967] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[968] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[969] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[970] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[971] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[972] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[973] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[974] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[975] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[976] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[977] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[978] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[979] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[980] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[981] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[982] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[983] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[984] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[985] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[986] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[987] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[988] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[989] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[990] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[991] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[992] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[993] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[994] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[995] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[996] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[997] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[998] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[999] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1000] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1001] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1002] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1003] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1004] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1005] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1006] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1007] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1008] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1009] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1010] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1011] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1012] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1013] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1014] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1015] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1016] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1017] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1018] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1019] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1020] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1021] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1022] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1023] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1024] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1025] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1026] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1027] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1028] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1029] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1030] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1031] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1032] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1033] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1034] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1035] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1036] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1037] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1038] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1039] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1040] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1041] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1042] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1043] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1044] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1045] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1046] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1047] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1048] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1049] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1050] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1051] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1052] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1053] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1054] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1055] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1056] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1057] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1058] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1059] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1060] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1061] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1062] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1063] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1064] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1065] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1066] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1067] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1068] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1069] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1070] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1071] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1072] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1073] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1074] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1075] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1076] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1077] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1078] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1079] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1080] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1081] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1082] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1083] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1084] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1085] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1086] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1087] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1088] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1089] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1090] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1091] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1092] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1093] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1094] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1095] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1096] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1097] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1098] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1099] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1100] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1101] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1102] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1103] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1104] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1105] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1106] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1107] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1108] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1109] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1110] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1111] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1112] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1113] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1114] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1115] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1116] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1117] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1118] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1119] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1120] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1121] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1122] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1123] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1124] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1125] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1126] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1127] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1128] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1129] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1130] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1131] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1132] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1133] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1134] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1135] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1136] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1137] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1138] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1139] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1140] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1141] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1142] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1143] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1144] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1145] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1146] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1147] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1148] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1149] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1150] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1151] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1152] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1153] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1154] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1155] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1156] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1157] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1158] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1159] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1160] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1161] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1162] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1163] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1164] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1165] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1166] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1167] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1168] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1169] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1170] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1171] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1172] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1173] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1174] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1175] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1176] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1177] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1178] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1179] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1180] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1181] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1182] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1183] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1184] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1185] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1186] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1187] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1188] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1189] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1190] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1191] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1192] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1193] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1194] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1195] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1196] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1197] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1198] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1199] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1200] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1201] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1202] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1203] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1204] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1205] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1206] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1207] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1208] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1209] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1210] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1211] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1212] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1213] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1214] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1215] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1216] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1217] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1218] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1219] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1220] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1221] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1222] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1223] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1224] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1225] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1226] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1227] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1228] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1229] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1230] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1231] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1232] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1233] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1234] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1235] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1236] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1237] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1238] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1239] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1240] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1241] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1242] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1243] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1244] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1245] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1246] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1247] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1248] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1249] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1250] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1251] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1252] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1253] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1254] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1255] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1256] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1257] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1258] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1259] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1260] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1261] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1262] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1263] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1264] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1265] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1266] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1267] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1268] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1269] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1270] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1271] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1272] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1273] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1274] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1275] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1276] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1277] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1278] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1279] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1280] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1281] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1282] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1283] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1284] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1285] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1286] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1287] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1288] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1289] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1290] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1291] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1292] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1293] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1294] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1295] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1296] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1297] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1298] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1299] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1300] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1301] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1302] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1303] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1304] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1305] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1306] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1307] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1308] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1309] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1310] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1311] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1312] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1313] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1314] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1315] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1316] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1317] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1318] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1319] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1320] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1321] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1322] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1323] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1324] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1325] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1326] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1327] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1328] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1329] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1330] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1331] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1332] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1333] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1334] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1335] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1336] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1337] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1338] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1339] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1340] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1341] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1342] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1343] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1344] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1345] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1346] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1347] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1348] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1349] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1350] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1351] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1352] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1353] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1354] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1355] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1356] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1357] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1358] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1359] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1360] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1361] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1362] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1363] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1364] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1365] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1366] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1367] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1368] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1369] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1370] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1371] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1372] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1373] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1374] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1375] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1376] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1377] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1378] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1379] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1380] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1381] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1382] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1383] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1384] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1385] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1386] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1387] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1388] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1389] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1390] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1391] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1392] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1393] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1394] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1395] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1396] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1397] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1398] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1399] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1400] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1401] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1402] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1403] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1404] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1405] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1406] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1407] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1408] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1409] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1410] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1411] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1412] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1413] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1414] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1415] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1416] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1417] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1418] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1419] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1420] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1421] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1422] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1423] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1424] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1425] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1426] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1427] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1428] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1429] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1430] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1431] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1432] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1433] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1434] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1435] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1436] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1437] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1438] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1439] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1440] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1441] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1442] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1443] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1444] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1445] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1446] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1447] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1448] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1449] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1450] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1451] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1452] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1453] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1454] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1455] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1456] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1457] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1458] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1459] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1460] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1461] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1462] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1463] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1464] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1465] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1466] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1467] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1468] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1469] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1470] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1471] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1472] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1473] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1474] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1475] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1476] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1477] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1478] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1479] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1480] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1481] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1482] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1483] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1484] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1485] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1486] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1487] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1488] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1489] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1490] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1491] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1492] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1493] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1494] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1495] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1496] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1497] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1498] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1499] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1500] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1501] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1502] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1503] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1504] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1505] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1506] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1507] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1508] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1509] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1510] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1511] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1512] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1513] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1514] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1515] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1516] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1517] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1518] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1519] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1520] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1521] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1522] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1523] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1524] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1525] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1526] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1527] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1528] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1529] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1530] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1531] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1532] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1533] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1534] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1535] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1536] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1537] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1538] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1539] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1540] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1541] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1542] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1543] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1544] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1545] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1546] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1547] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1548] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1549] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1550] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1551] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1552] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1553] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1554] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1555] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1556] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1557] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1558] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1559] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1560] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1561] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1562] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1563] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1564] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1565] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1566] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1567] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1568] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1569] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1570] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1571] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1572] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1573] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1574] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1575] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1576] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1577] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1578] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1579] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1580] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1581] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1582] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1583] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1584] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1585] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1586] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1587] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1588] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1589] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1590] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1591] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1592] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1593] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1594] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1595] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1596] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1597] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1598] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1599] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1600] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1601] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1602] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1603] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1604] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1605] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1606] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1607] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1608] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1609] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1610] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1611] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1612] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1613] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1614] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1615] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1616] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1617] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1618] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1619] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1620] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1621] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1622] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1623] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1624] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1625] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1626] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1627] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1628] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1629] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1630] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1631] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1632] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1633] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1634] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1635] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1636] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1637] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1638] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1639] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1640] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1641] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1642] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1643] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1644] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1645] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1646] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1647] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1648] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1649] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1650] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1651] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1652] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1653] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1654] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1655] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1656] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1657] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1658] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1659] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1660] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1661] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1662] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1663] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1664] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1665] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1666] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1667] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1668] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1669] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1670] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1671] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1672] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1673] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1674] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1675] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1676] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1677] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1678] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1679] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1680] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1681] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1682] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1683] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1684] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1685] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1686] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1687] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1688] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1689] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1690] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1691] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1692] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1693] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1694] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1695] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1696] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1697] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1698] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1699] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1700] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1701] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1702] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1703] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1704] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1705] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1706] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1707] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1708] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1709] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1710] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1711] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1712] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1713] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1714] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1715] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1716] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1717] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1718] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1719] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1720] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1721] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1722] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1723] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1724] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1725] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1726] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1727] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1728] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1729] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1730] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1731] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1732] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1733] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1734] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1735] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1736] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1737] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1738] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1739] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1740] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1741] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1742] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1743] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1744] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1745] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1746] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1747] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1748] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1749] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1750] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1751] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1752] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1753] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1754] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1755] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1756] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1757] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1758] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1759] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1760] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1761] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1762] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1763] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1764] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1765] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1766] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1767] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1768] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1769] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1770] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1771] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1772] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1773] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1774] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1775] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1776] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1777] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1778] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1779] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1780] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1781] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1782] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1783] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1784] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1785] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1786] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1787] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1788] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1789] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1790] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1791] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1792] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1793] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1794] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1795] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1796] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1797] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1798] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1799] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1800] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1801] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1802] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1803] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1804] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1805] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1806] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1807] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1808] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1809] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1810] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1811] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1812] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1813] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1814] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1815] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1816] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1817] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1818] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1819] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1820] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1821] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1822] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1823] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1824] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1825] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1826] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1827] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1828] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1829] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1830] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1831] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1832] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1833] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1834] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1835] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1836] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1837] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1838] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1839] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1840] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1841] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1842] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1843] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1844] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1845] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1846] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1847] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1848] = s[0] ? pos_SNs[17] : pos_SNs[17];
	assign level0[1849] = s[0] ? pos_SNs[17] : pos_SNs[17];
	assign level0[1850] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1851] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1852] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1853] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1854] = s[0] ? neg_SNs[22] : neg_SNs[22];
	assign level0[1855] = s[0] ? neg_SNs[22] : neg_SNs[22];
	assign level0[1856] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1857] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1858] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1859] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1860] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1861] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1862] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1863] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1864] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1865] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1866] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1867] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1868] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1869] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1870] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1871] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1872] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1873] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1874] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1875] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1876] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1877] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1878] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1879] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1880] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1881] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1882] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1883] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1884] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1885] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1886] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1887] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1888] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1889] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1890] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1891] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1892] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1893] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1894] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1895] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1896] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1897] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1898] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1899] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1900] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1901] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1902] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1903] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1904] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1905] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1906] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1907] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1908] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1909] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1910] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1911] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1912] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1913] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1914] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1915] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1916] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1917] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1918] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1919] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1920] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1921] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1922] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1923] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1924] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1925] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1926] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1927] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1928] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1929] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1930] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1931] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1932] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1933] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1934] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1935] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1936] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[1937] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[1938] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[1939] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[1940] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[1941] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[1942] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[1943] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[1944] = s[0] ? pos_SNs[131] : pos_SNs[131];
	assign level0[1945] = s[0] ? pos_SNs[131] : pos_SNs[131];
	assign level0[1946] = s[0] ? pos_SNs[14] : pos_SNs[14];
	assign level0[1947] = s[0] ? neg_SNs[15] : neg_SNs[15];
	assign level0[1948] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[1949] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1950] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1951] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1952] = s[0] ? neg_SNs[22] : neg_SNs[22];
	assign level0[1953] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1954] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1955] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1956] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1957] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1958] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1959] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1960] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1961] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1962] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[1963] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1964] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1965] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1966] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1967] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1968] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1969] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1970] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1971] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1972] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1973] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1974] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1975] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1976] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1977] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1978] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1979] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1980] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1981] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1982] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1983] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1984] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1985] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1986] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1987] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1988] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1989] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1990] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1991] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1992] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1993] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1994] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1995] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1996] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[1997] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[1998] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1999] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[2000] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[2001] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[2002] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[2003] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[2004] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[2005] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[2006] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[2007] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[2008] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2009] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[2010] = s[0] ? neg_SNs[132] : neg_SNs[132];
	assign level0[2011] = s[0] ? neg_SNs[133] : neg_SNs[133];
	assign level0[2012] = s[0] ? pos_SNs[134] : pos_SNs[134];
	assign level0[2013] = s[0] ? pos_SNs[10] : pos_SNs[10];
	assign level0[2014] = s[0] ? pos_SNs[13] : pos_SNs[13];
	assign level0[2015] = s[0] ? pos_SNs[17] : pos_SNs[17];
	assign level0[2016] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[2017] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[2018] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[2019] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[2020] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[2021] = s[0] ? neg_SNs[37] : neg_SNs[37];
	assign level0[2022] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[2023] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[2024] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[2025] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[2026] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[2027] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[2028] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[2029] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[2030] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[2031] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[2032] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[2033] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[2034] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[2035] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[2036] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[2037] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[2038] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[2039] = s[0] ? neg_SNs[110] : neg_SNs[110];
	assign level0[2040] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[2041] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[2042] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[2043] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[2044] = s[0] ? neg_SNs[126] : neg_SNs[126];
	assign level0[2045] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2046] = s[0] ? neg_SNs[133] : neg_SNs[133];
	assign level0[2047] = s[0] ? neg_SNs[136] : neg_SNs[136];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module hw_tree5  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[2] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[3] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[4] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[5] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[6] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[7] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[8] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[9] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[10] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[11] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[12] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[13] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[14] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[15] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[16] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[17] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[18] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[19] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[20] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[21] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[22] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[23] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[24] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[25] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[26] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[27] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[28] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[29] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[30] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[31] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[32] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[33] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[34] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[35] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[36] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[37] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[38] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[39] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[40] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[41] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[42] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[43] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[44] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[45] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[46] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[47] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[48] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[49] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[50] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[51] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[52] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[53] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[54] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[55] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[56] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[57] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[58] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[59] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[60] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[61] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[62] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[63] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[64] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[65] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[66] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[67] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[68] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[69] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[70] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[71] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[72] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[73] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[74] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[75] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[76] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[77] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[78] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[79] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[80] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[81] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[82] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[83] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[84] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[85] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[86] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[87] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[88] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[89] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[90] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[91] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[92] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[93] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[94] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[95] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[96] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[97] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[98] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[99] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[100] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[101] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[102] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[103] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[104] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[105] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[106] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[107] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[108] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[109] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[110] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[111] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[112] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[113] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[114] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[115] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[116] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[117] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[118] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[119] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[120] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[121] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[122] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[123] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[124] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[125] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[126] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[127] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[128] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[129] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[130] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[131] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[132] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[133] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[134] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[135] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[136] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[137] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[138] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[139] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[140] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[141] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[142] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[143] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[144] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[145] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[146] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[147] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[148] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[149] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[150] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[151] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[152] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[153] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[154] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[155] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[156] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[157] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[158] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[159] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[160] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[161] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[162] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[163] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[164] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[165] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[166] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[167] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[168] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[169] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[170] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[171] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[172] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[173] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[174] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[175] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[176] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[177] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[178] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[179] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[180] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[181] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[182] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[183] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[184] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[185] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[186] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[187] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[188] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[189] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[190] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[191] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[192] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[193] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[194] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[195] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[196] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[197] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[198] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[199] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[200] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[201] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[202] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[203] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[204] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[205] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[206] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[207] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[208] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[209] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[210] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[211] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[212] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[213] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[214] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[215] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[216] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[217] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[218] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[219] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[220] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[221] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[222] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[223] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[224] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[225] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[226] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[227] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[228] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[229] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[230] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[231] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[232] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[233] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[234] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[235] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[236] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[237] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[238] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[239] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[240] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[241] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[242] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[243] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[244] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[245] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[246] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[247] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[248] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[249] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[250] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[251] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[252] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[253] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[254] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[255] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[256] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[257] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[258] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[259] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[260] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[261] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[262] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[263] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[264] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[265] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[266] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[267] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[268] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[269] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[270] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[271] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[272] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[273] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[274] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[275] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[276] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[277] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[278] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[279] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[280] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[281] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[282] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[283] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[284] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[285] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[286] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[287] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[288] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[289] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[290] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[291] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[292] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[293] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[294] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[295] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[296] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[297] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[298] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[299] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[300] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[301] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[302] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[303] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[304] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[305] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[306] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[307] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[308] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[309] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[310] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[311] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[312] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[313] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[314] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[315] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[316] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[317] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[318] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[319] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[320] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[321] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[322] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[323] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[324] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[325] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[326] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[327] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[328] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[329] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[330] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[331] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[332] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[333] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[334] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[335] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[336] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[337] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[338] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[339] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[340] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[341] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[342] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[343] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[344] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[345] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[346] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[347] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[348] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[349] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[350] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[351] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[352] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[353] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[354] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[355] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[356] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[357] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[358] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[359] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[360] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[361] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[362] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[363] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[364] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[365] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[366] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[367] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[368] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[369] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[370] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[371] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[372] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[373] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[374] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[375] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[376] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[377] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[378] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[379] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[380] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[381] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[382] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[383] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[384] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[385] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[386] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[387] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[388] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[389] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[390] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[391] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[392] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[393] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[394] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[395] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[396] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[397] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[398] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[399] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[400] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[401] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[402] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[403] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[404] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[405] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[406] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[407] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[408] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[409] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[410] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[411] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[412] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[413] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[414] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[415] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[416] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[417] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[418] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[419] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[420] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[421] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[422] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[423] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[424] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[425] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[426] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[427] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[428] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[429] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[430] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[431] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[432] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[433] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[434] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[435] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[436] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[437] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[438] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[439] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[440] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[441] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[442] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[443] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[444] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[445] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[446] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[447] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[448] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[449] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[450] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[451] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[452] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[453] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[454] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[455] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[456] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[457] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[458] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[459] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[460] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[461] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[462] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[463] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[464] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[465] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[466] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[467] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[468] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[469] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[470] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[471] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[472] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[473] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[474] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[475] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[476] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[477] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[478] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[479] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[480] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[481] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[482] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[483] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[484] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[485] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[486] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[487] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[488] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[489] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[490] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[491] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[492] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[493] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[494] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[495] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[496] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[497] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[498] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[499] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[500] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[501] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[502] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[503] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[504] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[505] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[506] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[507] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[508] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[509] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[510] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[511] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[512] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[513] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[514] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[515] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[516] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[517] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[518] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[519] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[520] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[521] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[522] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[523] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[524] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[525] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[526] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[527] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[528] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[529] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[530] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[531] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[532] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[533] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[534] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[535] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[536] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[537] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[538] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[539] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[540] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[541] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[542] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[543] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[544] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[545] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[546] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[547] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[548] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[549] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[550] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[551] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[552] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[553] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[554] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[555] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[556] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[557] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[558] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[559] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[560] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[561] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[562] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[563] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[564] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[565] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[566] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[567] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[568] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[569] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[570] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[571] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[572] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[573] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[574] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[575] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[576] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[577] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[578] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[579] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[580] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[581] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[582] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[583] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[584] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[585] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[586] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[587] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[588] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[589] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[590] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[591] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[592] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[593] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[594] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[595] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[596] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[597] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[598] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[599] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[600] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[601] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[602] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[603] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[604] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[605] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[606] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[607] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[608] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[609] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[610] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[611] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[612] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[613] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[614] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[615] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[616] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[617] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[618] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[619] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[620] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[621] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[622] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[623] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[624] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[625] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[626] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[627] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[628] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[629] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[630] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[631] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[632] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[633] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[634] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[635] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[636] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[637] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[638] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[639] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[640] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[641] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[642] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[643] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[644] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[645] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[646] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[647] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[648] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[649] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[650] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[651] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[652] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[653] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[654] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[655] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[656] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[657] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[658] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[659] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[660] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[661] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[662] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[663] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[664] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[665] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[666] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[667] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[668] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[669] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[670] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[671] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[672] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[673] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[674] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[675] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[676] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[677] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[678] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[679] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[680] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[681] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[682] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[683] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[684] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[685] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[686] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[687] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[688] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[689] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[690] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[691] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[692] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[693] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[694] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[695] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[696] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[697] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[698] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[699] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[700] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[701] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[702] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[703] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[704] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[705] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[706] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[707] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[708] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[709] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[710] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[711] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[712] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[713] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[714] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[715] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[716] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[717] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[718] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[719] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[720] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[721] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[722] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[723] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[724] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[725] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[726] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[727] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[728] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[729] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[730] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[731] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[732] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[733] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[734] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[735] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[736] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[737] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[738] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[739] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[740] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[741] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[742] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[743] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[744] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[745] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[746] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[747] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[748] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[749] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[750] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[751] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[752] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[753] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[754] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[755] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[756] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[757] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[758] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[759] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[760] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[761] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[762] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[763] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[764] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[765] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[766] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[767] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[768] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[769] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[770] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[771] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[772] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[773] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[774] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[775] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[776] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[777] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[778] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[779] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[780] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[781] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[782] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[783] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[784] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[785] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[786] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[787] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[788] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[789] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[790] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[791] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[792] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[793] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[794] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[795] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[796] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[797] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[798] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[799] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[800] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[801] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[802] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[803] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[804] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[805] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[806] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[807] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[808] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[809] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[810] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[811] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[812] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[813] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[814] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[815] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[816] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[817] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[818] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[819] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[820] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[821] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[822] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[823] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[824] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[825] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[826] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[827] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[828] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[829] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[830] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[831] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[832] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[833] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[834] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[835] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[836] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[837] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[838] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[839] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[840] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[841] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[842] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[843] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[844] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[845] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[846] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[847] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[848] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[849] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[850] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[851] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[852] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[853] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[854] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[855] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[856] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[857] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[858] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[859] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[860] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[861] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[862] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[863] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[864] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[865] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[866] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[867] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[868] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[869] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[870] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[871] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[872] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[873] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[874] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[875] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[876] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[877] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[878] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[879] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[880] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[881] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[882] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[883] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[884] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[885] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[886] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[887] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[888] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[889] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[890] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[891] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[892] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[893] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[894] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[895] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[896] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[897] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[898] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[899] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[900] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[901] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[902] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[903] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[904] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[905] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[906] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[907] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[908] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[909] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[910] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[911] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[912] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[913] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[914] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[915] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[916] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[917] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[918] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[919] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[920] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[921] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[922] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[923] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[924] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[925] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[926] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[927] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[928] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[929] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[930] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[931] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[932] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[933] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[934] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[935] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[936] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[937] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[938] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[939] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[940] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[941] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[942] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[943] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[944] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[945] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[946] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[947] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[948] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[949] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[950] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[951] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[952] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[953] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[954] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[955] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[956] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[957] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[958] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[959] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[960] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[961] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[962] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[963] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[964] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[965] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[966] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[967] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[968] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[969] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[970] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[971] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[972] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[973] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[974] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[975] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[976] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[977] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[978] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[979] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[980] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[981] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[982] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[983] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[984] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[985] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[986] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[987] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[988] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[989] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[990] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[991] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[992] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[993] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[994] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[995] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[996] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[997] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[998] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[999] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1000] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1001] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1002] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1003] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1004] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1005] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1006] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1007] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1008] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1009] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1010] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1011] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1012] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1013] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1014] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1015] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1016] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1017] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1018] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1019] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1020] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1021] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1022] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1023] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1024] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1025] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1026] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1027] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1028] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1029] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1030] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1031] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1032] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1033] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1034] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1035] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1036] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1037] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1038] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1039] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1040] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1041] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1042] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1043] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1044] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1045] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1046] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1047] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1048] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1049] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1050] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1051] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1052] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1053] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1054] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1055] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1056] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1057] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1058] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1059] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1060] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1061] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1062] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1063] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1064] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1065] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1066] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1067] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1068] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1069] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1070] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1071] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1072] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1073] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1074] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1075] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1076] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1077] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1078] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1079] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1080] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1081] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1082] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1083] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1084] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1085] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1086] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1087] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1088] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1089] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1090] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1091] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1092] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1093] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1094] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1095] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1096] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1097] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1098] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1099] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1100] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1101] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1102] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1103] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1104] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1105] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1106] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1107] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1108] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1109] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1110] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1111] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1112] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1113] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1114] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1115] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1116] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1117] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1118] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1119] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1120] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1121] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1122] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1123] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1124] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1125] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1126] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1127] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1128] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1129] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1130] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1131] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1132] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1133] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1134] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1135] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1136] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1137] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1138] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1139] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1140] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1141] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1142] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1143] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1144] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1145] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1146] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1147] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1148] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1149] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1150] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1151] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1152] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1153] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1154] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1155] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1156] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1157] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1158] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1159] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1160] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1161] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1162] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1163] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1164] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1165] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1166] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1167] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1168] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1169] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1170] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1171] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1172] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1173] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1174] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1175] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1176] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1177] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1178] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1179] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1180] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1181] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1182] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1183] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1184] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1185] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1186] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1187] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1188] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1189] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1190] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1191] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1192] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1193] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1194] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1195] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1196] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1197] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1198] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1199] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1200] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1201] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1202] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1203] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1204] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1205] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1206] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1207] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1208] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1209] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1210] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1211] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1212] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1213] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1214] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1215] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1216] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1217] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1218] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1219] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1220] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1221] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1222] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1223] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1224] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1225] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1226] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1227] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1228] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1229] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1230] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1231] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1232] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1233] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1234] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1235] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1236] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1237] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1238] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1239] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1240] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1241] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1242] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1243] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1244] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1245] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1246] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1247] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1248] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1249] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1250] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1251] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1252] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1253] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1254] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1255] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1256] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1257] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1258] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1259] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1260] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1261] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1262] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1263] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1264] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1265] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1266] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1267] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1268] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1269] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1270] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1271] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1272] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1273] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1274] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1275] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1276] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1277] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1278] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1279] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1280] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1281] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1282] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1283] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1284] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1285] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1286] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1287] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1288] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1289] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1290] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1291] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1292] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1293] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1294] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1295] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1296] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1297] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1298] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1299] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1300] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1301] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1302] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1303] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1304] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1305] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1306] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1307] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1308] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1309] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1310] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1311] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1312] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1313] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1314] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1315] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1316] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1317] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1318] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1319] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1320] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1321] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1322] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1323] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1324] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1325] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1326] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1327] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1328] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1329] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1330] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1331] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1332] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1333] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1334] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1335] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1336] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1337] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1338] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1339] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1340] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1341] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1342] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1343] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1344] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1345] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1346] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1347] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1348] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1349] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1350] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1351] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1352] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1353] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1354] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1355] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1356] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1357] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1358] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1359] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1360] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1361] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1362] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1363] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1364] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1365] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1366] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1367] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1368] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1369] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1370] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1371] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1372] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1373] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1374] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1375] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1376] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1377] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1378] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1379] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1380] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1381] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1382] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1383] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1384] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1385] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1386] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1387] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1388] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1389] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1390] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1391] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1392] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1393] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1394] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1395] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1396] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1397] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1398] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1399] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1400] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1401] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1402] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1403] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1404] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1405] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1406] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1407] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1408] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1409] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1410] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1411] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1412] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1413] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1414] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1415] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1416] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1417] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1418] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1419] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1420] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1421] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1422] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1423] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1424] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1425] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1426] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1427] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1428] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1429] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1430] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1431] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1432] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1433] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1434] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1435] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1436] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1437] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1438] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1439] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1440] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1441] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1442] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1443] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1444] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1445] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1446] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1447] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1448] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1449] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1450] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1451] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1452] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1453] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1454] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1455] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1456] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1457] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1458] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1459] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1460] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1461] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1462] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1463] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1464] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1465] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1466] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1467] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1468] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1469] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1470] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1471] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1472] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1473] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1474] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1475] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1476] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1477] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1478] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1479] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1480] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1481] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1482] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1483] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1484] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1485] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1486] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1487] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1488] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1489] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1490] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1491] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1492] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1493] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1494] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1495] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1496] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1497] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1498] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1499] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1500] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1501] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1502] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1503] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1504] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1505] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1506] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1507] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1508] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1509] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1510] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1511] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1512] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1513] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1514] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1515] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1516] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1517] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1518] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1519] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1520] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1521] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1522] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1523] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1524] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1525] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1526] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1527] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1528] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1529] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1530] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1531] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1532] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1533] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1534] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1535] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1536] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1537] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1538] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1539] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1540] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1541] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1542] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1543] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1544] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1545] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1546] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1547] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1548] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1549] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1550] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1551] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1552] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1553] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1554] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1555] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1556] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1557] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1558] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1559] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1560] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1561] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1562] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1563] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1564] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1565] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1566] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1567] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1568] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1569] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1570] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1571] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1572] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1573] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1574] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1575] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1576] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1577] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1578] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1579] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1580] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1581] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1582] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1583] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1584] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1585] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1586] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1587] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1588] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1589] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1590] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1591] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1592] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1593] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1594] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1595] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1596] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1597] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1598] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1599] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1600] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1601] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1602] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1603] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1604] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1605] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1606] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1607] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1608] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1609] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1610] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1611] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1612] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1613] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1614] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1615] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1616] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1617] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1618] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1619] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1620] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1621] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1622] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1623] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1624] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1625] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1626] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1627] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1628] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1629] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1630] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1631] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1632] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1633] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1634] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1635] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1636] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1637] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1638] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1639] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1640] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1641] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1642] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1643] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1644] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1645] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1646] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1647] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1648] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1649] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1650] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1651] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1652] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1653] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1654] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1655] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1656] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1657] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1658] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1659] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1660] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1661] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1662] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1663] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1664] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1665] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1666] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1667] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1668] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1669] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1670] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1671] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1672] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1673] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1674] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1675] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1676] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1677] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1678] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1679] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1680] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1681] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1682] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1683] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1684] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1685] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1686] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1687] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1688] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1689] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1690] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1691] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1692] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1693] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1694] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1695] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1696] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1697] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1698] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1699] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1700] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1701] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1702] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1703] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1704] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1705] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1706] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1707] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1708] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1709] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1710] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1711] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1712] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1713] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1714] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1715] = s[0] ? pos_SNs[44] : pos_SNs[44];
	assign level0[1716] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1717] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1718] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1719] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1720] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1721] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1722] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1723] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1724] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1725] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1726] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1727] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1728] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1729] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1730] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1731] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1732] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1733] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1734] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1735] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1736] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1737] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1738] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1739] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1740] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1741] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1742] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1743] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1744] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1745] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1746] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1747] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1748] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1749] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1750] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1751] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1752] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1753] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1754] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1755] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1756] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1757] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1758] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1759] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1760] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1761] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1762] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1763] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1764] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1765] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1766] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1767] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1768] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1769] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1770] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1771] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1772] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1773] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1774] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1775] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1776] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1777] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1778] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1779] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1780] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1781] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1782] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1783] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1784] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1785] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1786] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1787] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1788] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1789] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1790] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1791] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1792] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1793] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1794] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1795] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1796] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1797] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1798] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1799] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1800] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1801] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1802] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1803] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1804] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1805] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1806] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1807] = s[0] ? pos_SNs[104] : pos_SNs[104];
	assign level0[1808] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1809] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1810] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1811] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1812] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1813] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1814] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1815] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1816] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1817] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1818] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1819] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[1820] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1821] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1822] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1823] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[1824] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1825] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1826] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1827] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1828] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1829] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1830] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1831] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1832] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1833] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1834] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1835] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1836] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1837] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1838] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1839] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1840] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1841] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1842] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1843] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1844] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[1845] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[1846] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[1847] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[1848] = s[0] ? pos_SNs[16] : pos_SNs[16];
	assign level0[1849] = s[0] ? pos_SNs[16] : pos_SNs[16];
	assign level0[1850] = s[0] ? neg_SNs[17] : neg_SNs[17];
	assign level0[1851] = s[0] ? neg_SNs[17] : neg_SNs[17];
	assign level0[1852] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1853] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1854] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[1855] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[1856] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1857] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1858] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1859] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1860] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1861] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1862] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1863] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1864] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1865] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1866] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1867] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1868] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1869] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1870] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1871] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1872] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1873] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1874] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1875] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1876] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1877] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1878] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1879] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1880] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1881] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1882] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1883] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1884] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1885] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1886] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1887] = s[0] ? pos_SNs[60] : pos_SNs[60];
	assign level0[1888] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1889] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1890] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1891] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1892] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1893] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1894] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1895] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1896] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1897] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1898] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1899] = s[0] ? neg_SNs[72] : neg_SNs[72];
	assign level0[1900] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1901] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1902] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1903] = s[0] ? neg_SNs[76] : neg_SNs[76];
	assign level0[1904] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1905] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1906] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1907] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1908] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1909] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1910] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1911] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1912] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1913] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1914] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1915] = s[0] ? pos_SNs[88] : pos_SNs[88];
	assign level0[1916] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1917] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1918] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1919] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1920] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1921] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1922] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1923] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1924] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1925] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1926] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1927] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1928] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1929] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1930] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1931] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1932] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1933] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1934] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1935] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1936] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1937] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[1938] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1939] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1940] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[1941] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[1942] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1943] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[1944] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1945] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1946] = s[0] ? neg_SNs[128] : neg_SNs[128];
	assign level0[1947] = s[0] ? neg_SNs[128] : neg_SNs[128];
	assign level0[1948] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[1949] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[1950] = s[0] ? neg_SNs[131] : neg_SNs[131];
	assign level0[1951] = s[0] ? neg_SNs[131] : neg_SNs[131];
	assign level0[1952] = s[0] ? pos_SNs[132] : pos_SNs[132];
	assign level0[1953] = s[0] ? pos_SNs[132] : pos_SNs[132];
	assign level0[1954] = s[0] ? pos_SNs[13] : pos_SNs[13];
	assign level0[1955] = s[0] ? neg_SNs[14] : neg_SNs[14];
	assign level0[1956] = s[0] ? pos_SNs[19] : pos_SNs[19];
	assign level0[1957] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[1958] = s[0] ? pos_SNs[21] : pos_SNs[21];
	assign level0[1959] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1960] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1961] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1962] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1963] = s[0] ? pos_SNs[28] : pos_SNs[28];
	assign level0[1964] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1965] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1966] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1967] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1968] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1969] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[1970] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1971] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1972] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1973] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1974] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1975] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1976] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1977] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1978] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1979] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1980] = s[0] ? neg_SNs[54] : neg_SNs[54];
	assign level0[1981] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1982] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1983] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1984] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1985] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1986] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1987] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1988] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1989] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1990] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1991] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1992] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1993] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1994] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1995] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1996] = s[0] ? neg_SNs[94] : neg_SNs[94];
	assign level0[1997] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1998] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1999] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[2000] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[2001] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[2002] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[2003] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[2004] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[2005] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[2006] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[2007] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[2008] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[2009] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[2010] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[2011] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[2012] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[2013] = s[0] ? pos_SNs[120] : pos_SNs[120];
	assign level0[2014] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[2015] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[2016] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[2017] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2018] = s[0] ? pos_SNs[127] : pos_SNs[127];
	assign level0[2019] = s[0] ? neg_SNs[128] : neg_SNs[128];
	assign level0[2020] = s[0] ? pos_SNs[129] : pos_SNs[129];
	assign level0[2021] = s[0] ? neg_SNs[134] : neg_SNs[134];
	assign level0[2022] = s[0] ? pos_SNs[135] : pos_SNs[135];
	assign level0[2023] = s[0] ? pos_SNs[10] : pos_SNs[10];
	assign level0[2024] = s[0] ? neg_SNs[12] : neg_SNs[12];
	assign level0[2025] = s[0] ? neg_SNs[20] : neg_SNs[20];
	assign level0[2026] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[2027] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[2028] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[2029] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[2030] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[2031] = s[0] ? neg_SNs[38] : neg_SNs[38];
	assign level0[2032] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[2033] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[2034] = s[0] ? neg_SNs[54] : neg_SNs[54];
	assign level0[2035] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[2036] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[2037] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[2038] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[2039] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[2040] = s[0] ? neg_SNs[111] : neg_SNs[111];
	assign level0[2041] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[2042] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[2043] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[2044] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[2045] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2046] = s[0] ? neg_SNs[133] : neg_SNs[133];
	assign level0[2047] = s[0] ? neg_SNs[137] : neg_SNs[137];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module hw_tree6  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[2] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[3] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[4] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[5] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[6] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[7] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[8] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[9] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[10] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[11] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[12] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[13] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[14] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[15] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[16] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[17] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[18] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[19] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[20] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[21] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[22] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[23] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[24] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[25] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[26] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[27] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[28] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[29] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[30] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[31] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[32] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[33] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[34] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[35] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[36] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[37] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[38] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[39] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[40] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[41] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[42] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[43] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[44] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[45] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[46] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[47] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[48] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[49] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[50] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[51] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[52] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[53] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[54] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[55] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[56] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[57] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[58] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[59] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[60] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[61] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[62] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[63] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[64] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[65] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[66] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[67] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[68] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[69] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[70] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[71] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[72] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[73] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[74] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[75] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[76] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[77] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[78] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[79] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[80] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[81] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[82] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[83] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[84] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[85] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[86] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[87] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[88] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[89] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[90] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[91] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[92] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[93] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[94] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[95] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[96] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[97] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[98] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[99] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[100] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[101] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[102] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[103] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[104] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[105] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[106] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[107] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[108] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[109] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[110] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[111] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[112] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[113] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[114] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[115] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[116] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[117] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[118] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[119] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[120] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[121] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[122] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[123] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[124] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[125] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[126] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[127] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[128] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[129] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[130] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[131] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[132] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[133] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[134] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[135] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[136] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[137] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[138] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[139] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[140] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[141] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[142] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[143] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[144] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[145] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[146] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[147] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[148] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[149] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[150] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[151] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[152] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[153] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[154] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[155] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[156] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[157] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[158] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[159] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[160] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[161] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[162] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[163] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[164] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[165] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[166] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[167] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[168] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[169] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[170] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[171] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[172] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[173] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[174] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[175] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[176] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[177] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[178] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[179] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[180] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[181] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[182] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[183] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[184] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[185] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[186] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[187] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[188] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[189] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[190] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[191] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[192] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[193] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[194] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[195] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[196] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[197] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[198] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[199] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[200] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[201] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[202] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[203] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[204] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[205] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[206] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[207] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[208] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[209] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[210] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[211] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[212] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[213] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[214] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[215] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[216] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[217] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[218] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[219] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[220] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[221] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[222] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[223] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[224] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[225] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[226] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[227] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[228] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[229] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[230] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[231] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[232] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[233] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[234] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[235] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[236] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[237] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[238] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[239] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[240] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[241] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[242] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[243] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[244] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[245] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[246] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[247] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[248] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[249] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[250] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[251] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[252] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[253] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[254] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[255] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[256] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[257] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[258] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[259] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[260] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[261] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[262] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[263] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[264] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[265] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[266] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[267] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[268] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[269] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[270] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[271] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[272] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[273] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[274] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[275] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[276] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[277] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[278] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[279] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[280] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[281] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[282] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[283] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[284] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[285] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[286] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[287] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[288] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[289] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[290] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[291] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[292] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[293] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[294] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[295] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[296] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[297] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[298] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[299] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[300] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[301] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[302] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[303] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[304] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[305] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[306] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[307] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[308] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[309] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[310] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[311] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[312] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[313] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[314] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[315] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[316] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[317] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[318] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[319] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[320] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[321] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[322] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[323] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[324] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[325] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[326] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[327] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[328] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[329] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[330] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[331] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[332] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[333] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[334] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[335] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[336] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[337] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[338] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[339] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[340] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[341] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[342] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[343] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[344] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[345] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[346] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[347] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[348] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[349] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[350] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[351] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[352] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[353] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[354] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[355] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[356] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[357] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[358] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[359] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[360] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[361] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[362] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[363] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[364] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[365] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[366] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[367] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[368] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[369] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[370] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[371] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[372] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[373] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[374] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[375] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[376] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[377] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[378] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[379] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[380] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[381] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[382] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[383] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[384] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[385] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[386] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[387] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[388] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[389] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[390] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[391] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[392] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[393] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[394] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[395] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[396] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[397] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[398] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[399] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[400] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[401] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[402] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[403] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[404] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[405] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[406] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[407] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[408] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[409] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[410] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[411] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[412] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[413] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[414] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[415] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[416] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[417] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[418] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[419] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[420] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[421] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[422] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[423] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[424] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[425] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[426] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[427] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[428] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[429] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[430] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[431] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[432] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[433] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[434] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[435] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[436] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[437] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[438] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[439] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[440] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[441] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[442] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[443] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[444] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[445] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[446] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[447] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[448] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[449] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[450] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[451] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[452] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[453] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[454] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[455] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[456] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[457] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[458] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[459] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[460] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[461] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[462] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[463] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[464] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[465] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[466] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[467] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[468] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[469] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[470] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[471] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[472] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[473] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[474] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[475] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[476] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[477] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[478] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[479] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[480] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[481] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[482] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[483] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[484] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[485] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[486] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[487] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[488] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[489] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[490] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[491] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[492] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[493] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[494] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[495] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[496] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[497] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[498] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[499] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[500] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[501] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[502] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[503] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[504] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[505] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[506] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[507] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[508] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[509] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[510] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[511] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[512] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[513] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[514] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[515] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[516] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[517] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[518] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[519] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[520] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[521] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[522] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[523] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[524] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[525] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[526] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[527] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[528] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[529] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[530] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[531] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[532] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[533] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[534] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[535] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[536] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[537] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[538] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[539] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[540] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[541] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[542] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[543] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[544] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[545] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[546] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[547] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[548] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[549] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[550] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[551] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[552] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[553] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[554] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[555] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[556] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[557] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[558] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[559] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[560] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[561] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[562] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[563] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[564] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[565] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[566] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[567] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[568] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[569] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[570] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[571] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[572] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[573] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[574] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[575] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[576] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[577] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[578] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[579] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[580] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[581] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[582] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[583] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[584] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[585] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[586] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[587] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[588] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[589] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[590] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[591] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[592] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[593] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[594] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[595] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[596] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[597] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[598] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[599] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[600] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[601] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[602] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[603] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[604] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[605] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[606] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[607] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[608] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[609] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[610] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[611] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[612] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[613] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[614] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[615] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[616] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[617] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[618] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[619] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[620] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[621] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[622] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[623] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[624] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[625] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[626] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[627] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[628] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[629] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[630] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[631] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[632] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[633] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[634] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[635] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[636] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[637] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[638] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[639] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[640] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[641] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[642] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[643] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[644] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[645] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[646] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[647] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[648] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[649] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[650] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[651] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[652] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[653] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[654] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[655] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[656] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[657] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[658] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[659] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[660] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[661] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[662] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[663] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[664] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[665] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[666] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[667] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[668] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[669] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[670] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[671] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[672] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[673] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[674] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[675] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[676] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[677] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[678] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[679] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[680] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[681] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[682] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[683] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[684] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[685] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[686] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[687] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[688] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[689] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[690] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[691] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[692] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[693] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[694] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[695] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[696] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[697] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[698] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[699] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[700] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[701] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[702] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[703] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[704] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[705] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[706] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[707] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[708] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[709] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[710] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[711] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[712] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[713] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[714] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[715] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[716] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[717] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[718] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[719] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[720] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[721] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[722] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[723] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[724] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[725] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[726] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[727] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[728] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[729] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[730] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[731] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[732] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[733] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[734] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[735] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[736] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[737] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[738] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[739] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[740] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[741] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[742] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[743] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[744] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[745] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[746] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[747] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[748] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[749] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[750] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[751] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[752] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[753] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[754] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[755] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[756] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[757] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[758] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[759] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[760] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[761] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[762] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[763] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[764] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[765] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[766] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[767] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[768] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[769] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[770] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[771] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[772] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[773] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[774] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[775] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[776] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[777] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[778] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[779] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[780] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[781] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[782] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[783] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[784] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[785] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[786] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[787] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[788] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[789] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[790] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[791] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[792] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[793] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[794] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[795] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[796] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[797] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[798] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[799] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[800] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[801] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[802] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[803] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[804] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[805] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[806] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[807] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[808] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[809] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[810] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[811] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[812] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[813] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[814] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[815] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[816] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[817] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[818] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[819] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[820] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[821] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[822] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[823] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[824] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[825] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[826] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[827] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[828] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[829] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[830] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[831] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[832] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[833] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[834] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[835] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[836] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[837] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[838] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[839] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[840] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[841] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[842] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[843] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[844] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[845] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[846] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[847] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[848] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[849] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[850] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[851] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[852] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[853] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[854] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[855] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[856] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[857] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[858] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[859] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[860] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[861] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[862] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[863] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[864] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[865] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[866] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[867] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[868] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[869] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[870] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[871] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[872] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[873] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[874] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[875] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[876] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[877] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[878] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[879] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[880] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[881] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[882] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[883] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[884] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[885] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[886] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[887] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[888] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[889] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[890] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[891] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[892] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[893] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[894] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[895] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[896] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[897] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[898] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[899] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[900] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[901] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[902] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[903] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[904] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[905] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[906] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[907] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[908] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[909] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[910] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[911] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[912] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[913] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[914] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[915] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[916] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[917] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[918] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[919] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[920] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[921] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[922] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[923] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[924] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[925] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[926] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[927] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[928] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[929] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[930] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[931] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[932] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[933] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[934] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[935] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[936] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[937] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[938] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[939] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[940] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[941] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[942] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[943] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[944] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[945] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[946] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[947] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[948] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[949] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[950] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[951] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[952] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[953] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[954] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[955] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[956] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[957] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[958] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[959] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[960] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[961] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[962] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[963] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[964] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[965] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[966] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[967] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[968] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[969] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[970] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[971] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[972] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[973] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[974] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[975] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[976] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[977] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[978] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[979] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[980] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[981] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[982] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[983] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[984] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[985] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[986] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[987] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[988] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[989] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[990] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[991] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[992] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[993] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[994] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[995] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[996] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[997] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[998] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[999] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1000] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1001] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1002] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1003] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1004] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1005] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1006] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1007] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1008] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1009] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1010] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1011] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1012] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1013] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1014] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1015] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1016] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1017] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1018] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1019] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1020] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1021] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1022] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1023] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1024] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1025] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1026] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1027] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1028] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1029] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1030] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1031] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1032] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1033] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1034] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1035] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1036] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1037] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1038] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1039] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1040] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1041] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1042] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1043] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1044] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1045] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1046] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1047] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1048] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1049] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1050] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1051] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1052] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1053] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1054] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1055] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1056] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1057] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1058] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1059] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1060] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1061] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1062] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1063] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1064] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1065] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1066] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1067] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1068] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1069] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1070] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1071] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1072] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1073] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1074] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1075] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1076] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1077] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1078] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1079] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1080] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1081] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1082] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1083] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1084] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1085] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1086] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1087] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1088] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1089] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1090] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1091] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1092] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1093] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1094] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1095] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1096] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1097] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1098] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1099] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1100] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1101] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1102] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1103] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1104] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1105] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1106] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1107] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1108] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1109] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1110] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1111] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1112] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1113] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1114] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1115] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1116] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1117] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1118] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1119] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1120] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1121] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1122] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1123] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1124] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1125] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1126] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1127] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1128] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1129] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1130] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1131] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1132] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1133] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1134] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1135] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1136] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1137] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1138] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1139] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1140] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1141] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1142] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1143] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1144] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1145] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1146] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1147] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1148] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1149] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1150] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1151] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1152] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1153] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1154] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1155] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1156] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1157] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1158] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1159] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1160] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1161] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1162] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1163] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1164] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1165] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1166] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1167] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1168] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1169] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1170] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1171] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1172] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1173] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1174] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1175] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1176] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1177] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1178] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1179] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1180] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1181] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1182] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1183] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1184] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1185] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1186] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1187] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1188] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1189] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1190] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1191] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1192] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1193] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1194] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1195] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1196] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1197] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1198] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1199] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1200] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1201] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1202] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1203] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1204] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1205] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1206] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1207] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1208] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1209] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1210] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1211] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1212] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1213] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1214] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1215] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1216] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1217] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1218] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1219] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1220] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1221] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1222] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1223] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1224] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1225] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1226] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1227] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1228] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1229] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1230] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1231] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1232] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1233] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1234] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1235] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1236] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1237] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1238] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1239] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1240] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1241] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1242] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1243] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1244] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1245] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1246] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1247] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1248] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1249] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1250] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1251] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1252] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1253] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1254] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1255] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1256] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1257] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1258] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1259] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1260] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1261] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1262] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1263] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1264] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1265] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1266] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1267] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1268] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1269] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1270] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1271] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1272] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1273] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1274] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1275] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1276] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1277] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1278] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1279] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1280] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1281] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1282] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1283] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1284] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1285] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1286] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1287] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1288] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1289] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1290] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1291] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1292] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1293] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1294] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1295] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1296] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1297] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1298] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1299] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1300] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1301] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1302] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1303] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1304] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1305] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1306] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1307] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1308] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1309] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1310] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1311] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1312] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1313] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1314] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1315] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1316] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1317] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1318] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1319] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1320] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1321] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1322] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1323] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1324] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1325] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1326] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1327] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1328] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1329] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1330] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1331] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1332] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1333] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1334] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1335] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1336] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1337] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1338] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1339] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1340] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1341] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1342] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1343] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1344] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1345] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1346] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1347] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1348] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1349] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1350] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1351] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1352] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1353] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1354] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1355] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1356] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1357] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1358] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1359] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1360] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1361] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1362] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1363] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1364] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1365] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1366] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1367] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1368] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1369] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1370] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1371] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1372] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1373] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1374] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1375] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1376] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1377] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1378] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1379] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1380] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1381] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1382] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1383] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1384] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1385] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1386] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1387] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1388] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1389] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1390] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1391] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1392] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1393] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1394] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1395] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1396] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1397] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1398] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1399] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1400] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1401] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1402] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1403] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1404] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1405] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1406] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1407] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1408] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1409] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1410] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1411] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1412] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1413] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1414] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1415] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1416] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1417] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1418] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1419] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1420] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1421] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1422] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1423] = s[0] ? neg_SNs[52] : neg_SNs[52];
	assign level0[1424] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1425] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1426] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1427] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1428] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1429] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1430] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1431] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1432] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1433] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1434] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1435] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1436] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1437] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1438] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1439] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1440] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1441] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1442] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1443] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1444] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1445] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1446] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1447] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1448] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1449] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1450] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1451] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1452] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1453] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1454] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1455] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1456] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1457] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1458] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1459] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1460] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1461] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1462] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1463] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1464] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1465] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1466] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1467] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1468] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1469] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1470] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1471] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1472] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1473] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1474] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1475] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1476] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1477] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1478] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1479] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1480] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1481] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1482] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1483] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1484] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1485] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1486] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1487] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1488] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1489] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1490] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1491] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1492] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1493] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1494] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1495] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1496] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1497] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1498] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1499] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1500] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1501] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1502] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1503] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1504] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1505] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1506] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1507] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1508] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1509] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1510] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1511] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1512] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1513] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1514] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1515] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1516] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1517] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1518] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1519] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1520] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1521] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1522] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1523] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1524] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1525] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1526] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1527] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1528] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1529] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1530] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1531] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1532] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1533] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1534] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1535] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1536] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1537] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1538] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1539] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1540] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1541] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1542] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1543] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1544] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1545] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1546] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1547] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1548] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1549] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1550] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1551] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1552] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1553] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1554] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1555] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1556] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1557] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1558] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1559] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1560] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1561] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1562] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1563] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1564] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1565] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1566] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1567] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1568] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1569] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1570] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1571] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1572] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1573] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1574] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1575] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1576] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1577] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1578] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1579] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1580] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1581] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1582] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1583] = s[0] ? neg_SNs[96] : neg_SNs[96];
	assign level0[1584] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1585] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1586] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1587] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1588] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1589] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1590] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1591] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1592] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1593] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1594] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1595] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1596] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1597] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1598] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1599] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1600] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1601] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1602] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1603] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1604] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1605] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1606] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1607] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[1608] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1609] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1610] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1611] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1612] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1613] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1614] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1615] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1616] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1617] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1618] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1619] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1620] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1621] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1622] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1623] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1624] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1625] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1626] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1627] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1628] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1629] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1630] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1631] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1632] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1633] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1634] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1635] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1636] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1637] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1638] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1639] = s[0] ? pos_SNs[41] : pos_SNs[41];
	assign level0[1640] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1641] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1642] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1643] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1644] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1645] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1646] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1647] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1648] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1649] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1650] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1651] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1652] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1653] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1654] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1655] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1656] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1657] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1658] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1659] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1660] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1661] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1662] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1663] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1664] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1665] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1666] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1667] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1668] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1669] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1670] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1671] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1672] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1673] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1674] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1675] = s[0] ? pos_SNs[57] : pos_SNs[57];
	assign level0[1676] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1677] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1678] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1679] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1680] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1681] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1682] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1683] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1684] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1685] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1686] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1687] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1688] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1689] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1690] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1691] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1692] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1693] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1694] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1695] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1696] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1697] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1698] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1699] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1700] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1701] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1702] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1703] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1704] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1705] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1706] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1707] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1708] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1709] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1710] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1711] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1712] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1713] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1714] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1715] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1716] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1717] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1718] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1719] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1720] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1721] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1722] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1723] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1724] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1725] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1726] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1727] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1728] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1729] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1730] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1731] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1732] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1733] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1734] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1735] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1736] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1737] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1738] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1739] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1740] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1741] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1742] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1743] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1744] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1745] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1746] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1747] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1748] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1749] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1750] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1751] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1752] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1753] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1754] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1755] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1756] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1757] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1758] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1759] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1760] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1761] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1762] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1763] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1764] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1765] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1766] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1767] = s[0] ? pos_SNs[91] : pos_SNs[91];
	assign level0[1768] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1769] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1770] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1771] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1772] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1773] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1774] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1775] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1776] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1777] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1778] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1779] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1780] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1781] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1782] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1783] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1784] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1785] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1786] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1787] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[1788] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1789] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1790] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1791] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1792] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1793] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1794] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1795] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1796] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1797] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1798] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1799] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1800] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1801] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1802] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1803] = s[0] ? pos_SNs[107] : pos_SNs[107];
	assign level0[1804] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1805] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1806] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1807] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1808] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1809] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1810] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1811] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1812] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1813] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1814] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1815] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1816] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1817] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1818] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1819] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1820] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1821] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1822] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1823] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1824] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[1825] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[1826] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[1827] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[1828] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[1829] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[1830] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[1831] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[1832] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[1833] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[1834] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1835] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[1836] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1837] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1838] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1839] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1840] = s[0] ? neg_SNs[24] : neg_SNs[24];
	assign level0[1841] = s[0] ? neg_SNs[24] : neg_SNs[24];
	assign level0[1842] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1843] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1844] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1845] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1846] = s[0] ? neg_SNs[28] : neg_SNs[28];
	assign level0[1847] = s[0] ? neg_SNs[28] : neg_SNs[28];
	assign level0[1848] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1849] = s[0] ? neg_SNs[29] : neg_SNs[29];
	assign level0[1850] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1851] = s[0] ? pos_SNs[30] : pos_SNs[30];
	assign level0[1852] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1853] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1854] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1855] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[1856] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1857] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1858] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1859] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1860] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1861] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1862] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[1863] = s[0] ? pos_SNs[37] : pos_SNs[37];
	assign level0[1864] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1865] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1866] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1867] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1868] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1869] = s[0] ? neg_SNs[45] : neg_SNs[45];
	assign level0[1870] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1871] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1872] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1873] = s[0] ? pos_SNs[51] : pos_SNs[51];
	assign level0[1874] = s[0] ? neg_SNs[56] : neg_SNs[56];
	assign level0[1875] = s[0] ? neg_SNs[56] : neg_SNs[56];
	assign level0[1876] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1877] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1878] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1879] = s[0] ? pos_SNs[62] : pos_SNs[62];
	assign level0[1880] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1881] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1882] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1883] = s[0] ? neg_SNs[68] : neg_SNs[68];
	assign level0[1884] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1885] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1886] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1887] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[1888] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1889] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1890] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1891] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1892] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1893] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1894] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1895] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[1896] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1897] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1898] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1899] = s[0] ? neg_SNs[80] : neg_SNs[80];
	assign level0[1900] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1901] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1902] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1903] = s[0] ? pos_SNs[86] : pos_SNs[86];
	assign level0[1904] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1905] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1906] = s[0] ? neg_SNs[92] : neg_SNs[92];
	assign level0[1907] = s[0] ? neg_SNs[92] : neg_SNs[92];
	assign level0[1908] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1909] = s[0] ? pos_SNs[97] : pos_SNs[97];
	assign level0[1910] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1911] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1912] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1913] = s[0] ? neg_SNs[103] : neg_SNs[103];
	assign level0[1914] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1915] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1916] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1917] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[1918] = s[0] ? pos_SNs[111] : pos_SNs[111];
	assign level0[1919] = s[0] ? pos_SNs[111] : pos_SNs[111];
	assign level0[1920] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[1921] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[1922] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1923] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[1924] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1925] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[1926] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1927] = s[0] ? pos_SNs[116] : pos_SNs[116];
	assign level0[1928] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1929] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[1930] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1931] = s[0] ? pos_SNs[118] : pos_SNs[118];
	assign level0[1932] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1933] = s[0] ? neg_SNs[119] : neg_SNs[119];
	assign level0[1934] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[1935] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[1936] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1937] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[1938] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1939] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[1940] = s[0] ? neg_SNs[124] : neg_SNs[124];
	assign level0[1941] = s[0] ? neg_SNs[124] : neg_SNs[124];
	assign level0[1942] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1943] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[1944] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[1945] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[1946] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[1947] = s[0] ? neg_SNs[129] : neg_SNs[129];
	assign level0[1948] = s[0] ? neg_SNs[132] : neg_SNs[132];
	assign level0[1949] = s[0] ? neg_SNs[132] : neg_SNs[132];
	assign level0[1950] = s[0] ? neg_SNs[14] : neg_SNs[14];
	assign level0[1951] = s[0] ? pos_SNs[15] : pos_SNs[15];
	assign level0[1952] = s[0] ? pos_SNs[17] : pos_SNs[17];
	assign level0[1953] = s[0] ? pos_SNs[20] : pos_SNs[20];
	assign level0[1954] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1955] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1956] = s[0] ? pos_SNs[25] : pos_SNs[25];
	assign level0[1957] = s[0] ? neg_SNs[26] : neg_SNs[26];
	assign level0[1958] = s[0] ? neg_SNs[31] : neg_SNs[31];
	assign level0[1959] = s[0] ? neg_SNs[33] : neg_SNs[33];
	assign level0[1960] = s[0] ? pos_SNs[35] : pos_SNs[35];
	assign level0[1961] = s[0] ? neg_SNs[36] : neg_SNs[36];
	assign level0[1962] = s[0] ? neg_SNs[40] : neg_SNs[40];
	assign level0[1963] = s[0] ? neg_SNs[42] : neg_SNs[42];
	assign level0[1964] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1965] = s[0] ? pos_SNs[46] : pos_SNs[46];
	assign level0[1966] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[1967] = s[0] ? pos_SNs[48] : pos_SNs[48];
	assign level0[1968] = s[0] ? neg_SNs[49] : neg_SNs[49];
	assign level0[1969] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[1970] = s[0] ? neg_SNs[54] : neg_SNs[54];
	assign level0[1971] = s[0] ? neg_SNs[56] : neg_SNs[56];
	assign level0[1972] = s[0] ? neg_SNs[58] : neg_SNs[58];
	assign level0[1973] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1974] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1975] = s[0] ? neg_SNs[61] : neg_SNs[61];
	assign level0[1976] = s[0] ? neg_SNs[63] : neg_SNs[63];
	assign level0[1977] = s[0] ? pos_SNs[64] : pos_SNs[64];
	assign level0[1978] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[1979] = s[0] ? pos_SNs[67] : pos_SNs[67];
	assign level0[1980] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[1981] = s[0] ? neg_SNs[70] : neg_SNs[70];
	assign level0[1982] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1983] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1984] = s[0] ? neg_SNs[78] : neg_SNs[78];
	assign level0[1985] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[1986] = s[0] ? pos_SNs[81] : pos_SNs[81];
	assign level0[1987] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[1988] = s[0] ? pos_SNs[84] : pos_SNs[84];
	assign level0[1989] = s[0] ? neg_SNs[85] : neg_SNs[85];
	assign level0[1990] = s[0] ? neg_SNs[87] : neg_SNs[87];
	assign level0[1991] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1992] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1993] = s[0] ? neg_SNs[90] : neg_SNs[90];
	assign level0[1994] = s[0] ? neg_SNs[92] : neg_SNs[92];
	assign level0[1995] = s[0] ? neg_SNs[94] : neg_SNs[94];
	assign level0[1996] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[1997] = s[0] ? neg_SNs[99] : neg_SNs[99];
	assign level0[1998] = s[0] ? pos_SNs[100] : pos_SNs[100];
	assign level0[1999] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[2000] = s[0] ? pos_SNs[102] : pos_SNs[102];
	assign level0[2001] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[2002] = s[0] ? neg_SNs[106] : neg_SNs[106];
	assign level0[2003] = s[0] ? neg_SNs[108] : neg_SNs[108];
	assign level0[2004] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[2005] = s[0] ? pos_SNs[113] : pos_SNs[113];
	assign level0[2006] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[2007] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[2008] = s[0] ? neg_SNs[122] : neg_SNs[122];
	assign level0[2009] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[2010] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[2011] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2012] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2013] = s[0] ? pos_SNs[131] : pos_SNs[131];
	assign level0[2014] = s[0] ? pos_SNs[133] : pos_SNs[133];
	assign level0[2015] = s[0] ? neg_SNs[134] : neg_SNs[134];
	assign level0[2016] = s[0] ? neg_SNs[9] : neg_SNs[9];
	assign level0[2017] = s[0] ? neg_SNs[11] : neg_SNs[11];
	assign level0[2018] = s[0] ? pos_SNs[15] : pos_SNs[15];
	assign level0[2019] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[2020] = s[0] ? neg_SNs[24] : neg_SNs[24];
	assign level0[2021] = s[0] ? neg_SNs[28] : neg_SNs[28];
	assign level0[2022] = s[0] ? pos_SNs[32] : pos_SNs[32];
	assign level0[2023] = s[0] ? neg_SNs[34] : neg_SNs[34];
	assign level0[2024] = s[0] ? neg_SNs[38] : neg_SNs[38];
	assign level0[2025] = s[0] ? neg_SNs[47] : neg_SNs[47];
	assign level0[2026] = s[0] ? pos_SNs[53] : pos_SNs[53];
	assign level0[2027] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[2028] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[2029] = s[0] ? neg_SNs[65] : neg_SNs[65];
	assign level0[2030] = s[0] ? pos_SNs[69] : pos_SNs[69];
	assign level0[2031] = s[0] ? pos_SNs[71] : pos_SNs[71];
	assign level0[2032] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[2033] = s[0] ? pos_SNs[77] : pos_SNs[77];
	assign level0[2034] = s[0] ? pos_SNs[79] : pos_SNs[79];
	assign level0[2035] = s[0] ? neg_SNs[83] : neg_SNs[83];
	assign level0[2036] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[2037] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[2038] = s[0] ? pos_SNs[95] : pos_SNs[95];
	assign level0[2039] = s[0] ? neg_SNs[101] : neg_SNs[101];
	assign level0[2040] = s[0] ? neg_SNs[112] : neg_SNs[112];
	assign level0[2041] = s[0] ? neg_SNs[115] : neg_SNs[115];
	assign level0[2042] = s[0] ? neg_SNs[117] : neg_SNs[117];
	assign level0[2043] = s[0] ? pos_SNs[123] : pos_SNs[123];
	assign level0[2044] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2045] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2046] = s[0] ? pos_SNs[135] : pos_SNs[135];
	assign level0[2047] = s[0] ? pos_SNs[138] : pos_SNs[138];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module hw_tree7  (
	input  logic           pos_SNs  [148:0],
	input  logic           neg_SNs  [148:0],
	input  logic [11:0]     s,
	output logic           out
);
	logic level0  [2047:0];
	logic level1  [1023:0];
	logic level2  [511:0];
	logic level3  [255:0];
	logic level4  [127:0];
	logic level5  [63:0];
	logic level6  [31:0];
	logic level7  [15:0];
	logic level8  [7:0];
	logic level9  [3:0];
	logic level10  [1:0];
	logic level11  [0:0];

	assign level0[0] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[2] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[3] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[4] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[5] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[6] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[7] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[8] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[9] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[10] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[11] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[12] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[13] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[14] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[15] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[16] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[17] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[18] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[19] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[20] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[21] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[22] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[23] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[24] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[25] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[26] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[27] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[28] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[29] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[30] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[31] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[32] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[33] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[34] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[35] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[36] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[37] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[38] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[39] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[40] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[41] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[42] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[43] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[44] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[45] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[46] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[47] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[48] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[49] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[50] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[51] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[52] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[53] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[54] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[55] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[56] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[57] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[58] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[59] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[60] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[61] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[62] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[63] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[64] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[65] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[66] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[67] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[68] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[69] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[70] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[71] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[72] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[73] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[74] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[75] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[76] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[77] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[78] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[79] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[80] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[81] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[82] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[83] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[84] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[85] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[86] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[87] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[88] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[89] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[90] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[91] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[92] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[93] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[94] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[95] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[96] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[97] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[98] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[99] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[100] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[101] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[102] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[103] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[104] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[105] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[106] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[107] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[108] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[109] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[110] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[111] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[112] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[113] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[114] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[115] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[116] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[117] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[118] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[119] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[120] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[121] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[122] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[123] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[124] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[125] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[126] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[127] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[128] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[129] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[130] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[131] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[132] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[133] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[134] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[135] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[136] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[137] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[138] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[139] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[140] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[141] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[142] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[143] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[144] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[145] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[146] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[147] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[148] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[149] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[150] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[151] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[152] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[153] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[154] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[155] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[156] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[157] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[158] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[159] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[160] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[161] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[162] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[163] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[164] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[165] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[166] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[167] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[168] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[169] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[170] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[171] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[172] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[173] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[174] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[175] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[176] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[177] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[178] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[179] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[180] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[181] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[182] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[183] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[184] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[185] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[186] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[187] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[188] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[189] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[190] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[191] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[192] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[193] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[194] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[195] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[196] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[197] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[198] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[199] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[200] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[201] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[202] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[203] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[204] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[205] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[206] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[207] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[208] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[209] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[210] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[211] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[212] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[213] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[214] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[215] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[216] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[217] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[218] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[219] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[220] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[221] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[222] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[223] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[224] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[225] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[226] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[227] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[228] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[229] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[230] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[231] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[232] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[233] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[234] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[235] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[236] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[237] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[238] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[239] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[240] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[241] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[242] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[243] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[244] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[245] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[246] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[247] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[248] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[249] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[250] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[251] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[252] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[253] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[254] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[255] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[256] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[257] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[258] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[259] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[260] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[261] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[262] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[263] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[264] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[265] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[266] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[267] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[268] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[269] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[270] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[271] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[272] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[273] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[274] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[275] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[276] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[277] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[278] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[279] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[280] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[281] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[282] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[283] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[284] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[285] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[286] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[287] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[288] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[289] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[290] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[291] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[292] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[293] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[294] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[295] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[296] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[297] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[298] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[299] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[300] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[301] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[302] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[303] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[304] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[305] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[306] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[307] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[308] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[309] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[310] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[311] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[312] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[313] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[314] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[315] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[316] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[317] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[318] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[319] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[320] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[321] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[322] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[323] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[324] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[325] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[326] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[327] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[328] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[329] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[330] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[331] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[332] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[333] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[334] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[335] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[336] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[337] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[338] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[339] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[340] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[341] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[342] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[343] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[344] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[345] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[346] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[347] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[348] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[349] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[350] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[351] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[352] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[353] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[354] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[355] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[356] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[357] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[358] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[359] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[360] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[361] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[362] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[363] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[364] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[365] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[366] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[367] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[368] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[369] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[370] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[371] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[372] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[373] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[374] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[375] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[376] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[377] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[378] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[379] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[380] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[381] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[382] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[383] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[384] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[385] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[386] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[387] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[388] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[389] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[390] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[391] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[392] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[393] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[394] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[395] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[396] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[397] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[398] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[399] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[400] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[401] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[402] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[403] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[404] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[405] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[406] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[407] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[408] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[409] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[410] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[411] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[412] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[413] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[414] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[415] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[416] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[417] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[418] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[419] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[420] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[421] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[422] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[423] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[424] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[425] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[426] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[427] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[428] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[429] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[430] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[431] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[432] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[433] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[434] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[435] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[436] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[437] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[438] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[439] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[440] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[441] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[442] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[443] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[444] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[445] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[446] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[447] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[448] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[449] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[450] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[451] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[452] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[453] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[454] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[455] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[456] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[457] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[458] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[459] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[460] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[461] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[462] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[463] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[464] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[465] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[466] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[467] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[468] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[469] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[470] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[471] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[472] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[473] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[474] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[475] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[476] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[477] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[478] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[479] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[480] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[481] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[482] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[483] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[484] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[485] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[486] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[487] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[488] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[489] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[490] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[491] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[492] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[493] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[494] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[495] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[496] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[497] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[498] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[499] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[500] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[501] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[502] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[503] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[504] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[505] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[506] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[507] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[508] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[509] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[510] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[511] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[512] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[513] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[514] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[515] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[516] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[517] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[518] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[519] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[520] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[521] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[522] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[523] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[524] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[525] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[526] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[527] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[528] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[529] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[530] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[531] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[532] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[533] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[534] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[535] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[536] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[537] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[538] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[539] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[540] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[541] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[542] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[543] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[544] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[545] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[546] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[547] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[548] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[549] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[550] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[551] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[552] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[553] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[554] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[555] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[556] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[557] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[558] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[559] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[560] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[561] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[562] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[563] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[564] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[565] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[566] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[567] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[568] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[569] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[570] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[571] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[572] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[573] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[574] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[575] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[576] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[577] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[578] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[579] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[580] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[581] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[582] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[583] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[584] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[585] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[586] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[587] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[588] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[589] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[590] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[591] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[592] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[593] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[594] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[595] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[596] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[597] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[598] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[599] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[600] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[601] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[602] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[603] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[604] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[605] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[606] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[607] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[608] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[609] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[610] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[611] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[612] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[613] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[614] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[615] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[616] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[617] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[618] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[619] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[620] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[621] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[622] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[623] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[624] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[625] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[626] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[627] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[628] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[629] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[630] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[631] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[632] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[633] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[634] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[635] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[636] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[637] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[638] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[639] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[640] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[641] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[642] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[643] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[644] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[645] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[646] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[647] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[648] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[649] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[650] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[651] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[652] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[653] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[654] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[655] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[656] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[657] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[658] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[659] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[660] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[661] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[662] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[663] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[664] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[665] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[666] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[667] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[668] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[669] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[670] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[671] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[672] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[673] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[674] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[675] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[676] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[677] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[678] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[679] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[680] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[681] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[682] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[683] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[684] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[685] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[686] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[687] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[688] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[689] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[690] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[691] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[692] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[693] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[694] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[695] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[696] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[697] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[698] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[699] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[700] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[701] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[702] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[703] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[704] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[705] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[706] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[707] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[708] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[709] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[710] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[711] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[712] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[713] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[714] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[715] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[716] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[717] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[718] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[719] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[720] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[721] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[722] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[723] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[724] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[725] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[726] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[727] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[728] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[729] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[730] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[731] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[732] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[733] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[734] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[735] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[736] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[737] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[738] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[739] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[740] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[741] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[742] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[743] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[744] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[745] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[746] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[747] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[748] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[749] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[750] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[751] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[752] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[753] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[754] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[755] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[756] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[757] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[758] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[759] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[760] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[761] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[762] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[763] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[764] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[765] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[766] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[767] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[768] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[769] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[770] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[771] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[772] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[773] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[774] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[775] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[776] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[777] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[778] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[779] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[780] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[781] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[782] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[783] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[784] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[785] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[786] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[787] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[788] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[789] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[790] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[791] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[792] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[793] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[794] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[795] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[796] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[797] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[798] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[799] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[800] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[801] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[802] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[803] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[804] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[805] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[806] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[807] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[808] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[809] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[810] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[811] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[812] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[813] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[814] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[815] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[816] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[817] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[818] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[819] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[820] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[821] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[822] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[823] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[824] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[825] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[826] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[827] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[828] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[829] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[830] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[831] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[832] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[833] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[834] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[835] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[836] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[837] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[838] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[839] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[840] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[841] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[842] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[843] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[844] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[845] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[846] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[847] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[848] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[849] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[850] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[851] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[852] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[853] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[854] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[855] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[856] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[857] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[858] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[859] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[860] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[861] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[862] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[863] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[864] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[865] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[866] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[867] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[868] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[869] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[870] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[871] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[872] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[873] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[874] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[875] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[876] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[877] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[878] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[879] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[880] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[881] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[882] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[883] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[884] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[885] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[886] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[887] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[888] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[889] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[890] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[891] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[892] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[893] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[894] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[895] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[896] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[897] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[898] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[899] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[900] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[901] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[902] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[903] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[904] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[905] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[906] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[907] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[908] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[909] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[910] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[911] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[912] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[913] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[914] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[915] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[916] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[917] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[918] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[919] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[920] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[921] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[922] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[923] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[924] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[925] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[926] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[927] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[928] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[929] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[930] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[931] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[932] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[933] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[934] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[935] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[936] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[937] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[938] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[939] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[940] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[941] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[942] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[943] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[944] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[945] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[946] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[947] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[948] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[949] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[950] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[951] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[952] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[953] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[954] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[955] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[956] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[957] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[958] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[959] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[960] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[961] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[962] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[963] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[964] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[965] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[966] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[967] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[968] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[969] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[970] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[971] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[972] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[973] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[974] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[975] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[976] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[977] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[978] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[979] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[980] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[981] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[982] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[983] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[984] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[985] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[986] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[987] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[988] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[989] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[990] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[991] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[992] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[993] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[994] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[995] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[996] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[997] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[998] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[999] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1000] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1001] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1002] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1003] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1004] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1005] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1006] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1007] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1008] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1009] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1010] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1011] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1012] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1013] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1014] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1015] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1016] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1017] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1018] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1019] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1020] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1021] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1022] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1023] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1024] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1025] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1026] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1027] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1028] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1029] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1030] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1031] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1032] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1033] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1034] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1035] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1036] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1037] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1038] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1039] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1040] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1041] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1042] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1043] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1044] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1045] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1046] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1047] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1048] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1049] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1050] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1051] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1052] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1053] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1054] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1055] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1056] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1057] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1058] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1059] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1060] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1061] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1062] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1063] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1064] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1065] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1066] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1067] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1068] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1069] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1070] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1071] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1072] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1073] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1074] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1075] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1076] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1077] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1078] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1079] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1080] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1081] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1082] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1083] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1084] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1085] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1086] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1087] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1088] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1089] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1090] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1091] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1092] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1093] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1094] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1095] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1096] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1097] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1098] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1099] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1100] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1101] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1102] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1103] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1104] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1105] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1106] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1107] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1108] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1109] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1110] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1111] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1112] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1113] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1114] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1115] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1116] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1117] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1118] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1119] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1120] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1121] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1122] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1123] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1124] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1125] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1126] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1127] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1128] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1129] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1130] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1131] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1132] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1133] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1134] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1135] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1136] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1137] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1138] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1139] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1140] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1141] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1142] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1143] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1144] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1145] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1146] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1147] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1148] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1149] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1150] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1151] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1152] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1153] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1154] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1155] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1156] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1157] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1158] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1159] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1160] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1161] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1162] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1163] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1164] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1165] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1166] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1167] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1168] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1169] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1170] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1171] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1172] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1173] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1174] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1175] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1176] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1177] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1178] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1179] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1180] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1181] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1182] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1183] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1184] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1185] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1186] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1187] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1188] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1189] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1190] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1191] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1192] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1193] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1194] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1195] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1196] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1197] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1198] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1199] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1200] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1201] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1202] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1203] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1204] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1205] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1206] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1207] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1208] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1209] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1210] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1211] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1212] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1213] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1214] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1215] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1216] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1217] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1218] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1219] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1220] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1221] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1222] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1223] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1224] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1225] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1226] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1227] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1228] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1229] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1230] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1231] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1232] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1233] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1234] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1235] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1236] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1237] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1238] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1239] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1240] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1241] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1242] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1243] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1244] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1245] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1246] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1247] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1248] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1249] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1250] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1251] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1252] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1253] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1254] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1255] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1256] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1257] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1258] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1259] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1260] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1261] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1262] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1263] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1264] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1265] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1266] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1267] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1268] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1269] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1270] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1271] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1272] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1273] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1274] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1275] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1276] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1277] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1278] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1279] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1280] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1281] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1282] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1283] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1284] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1285] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1286] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1287] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1288] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1289] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1290] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1291] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1292] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1293] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1294] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1295] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1296] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1297] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1298] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1299] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1300] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1301] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1302] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1303] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1304] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1305] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1306] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1307] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1308] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1309] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1310] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1311] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1312] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1313] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1314] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1315] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1316] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1317] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1318] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1319] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1320] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1321] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1322] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1323] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1324] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1325] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1326] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1327] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1328] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1329] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1330] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1331] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1332] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1333] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1334] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1335] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1336] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1337] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1338] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1339] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1340] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1341] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1342] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1343] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1344] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1345] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1346] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1347] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1348] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1349] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1350] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1351] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1352] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1353] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1354] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1355] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1356] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1357] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1358] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1359] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1360] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1361] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1362] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1363] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1364] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1365] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1366] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1367] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1368] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1369] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1370] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1371] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1372] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1373] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1374] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1375] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1376] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1377] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1378] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1379] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1380] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1381] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1382] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1383] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1384] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1385] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1386] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1387] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1388] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1389] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1390] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1391] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1392] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1393] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1394] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1395] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1396] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1397] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1398] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1399] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1400] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1401] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1402] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1403] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1404] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1405] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1406] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1407] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1408] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1409] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1410] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1411] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1412] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1413] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1414] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1415] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1416] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1417] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1418] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1419] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1420] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1421] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1422] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1423] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1424] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1425] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1426] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1427] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1428] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1429] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1430] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1431] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1432] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1433] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1434] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1435] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1436] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1437] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1438] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1439] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1440] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1441] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1442] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1443] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1444] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1445] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1446] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1447] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1448] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1449] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1450] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1451] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1452] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1453] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1454] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1455] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1456] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1457] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1458] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1459] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1460] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1461] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1462] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1463] = s[0] ? neg_SNs[46] : neg_SNs[46];
	assign level0[1464] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1465] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1466] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1467] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1468] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1469] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1470] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1471] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[1472] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1473] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1474] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1475] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1476] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1477] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1478] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1479] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1480] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1481] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1482] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1483] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1484] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1485] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1486] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1487] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1488] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1489] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1490] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1491] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1492] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1493] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1494] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1495] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1496] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1497] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1498] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1499] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1500] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1501] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1502] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1503] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1504] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1505] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1506] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1507] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1508] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1509] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1510] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1511] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1512] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1513] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1514] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1515] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1516] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1517] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1518] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1519] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[1520] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1521] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1522] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1523] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1524] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1525] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1526] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1527] = s[0] ? pos_SNs[61] : pos_SNs[61];
	assign level0[1528] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1529] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1530] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1531] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1532] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1533] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1534] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1535] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1536] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1537] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1538] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1539] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1540] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1541] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1542] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1543] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1544] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1545] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1546] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1547] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1548] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1549] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1550] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1551] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1552] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1553] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1554] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1555] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1556] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1557] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1558] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1559] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1560] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1561] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1562] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1563] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1564] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1565] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1566] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1567] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1568] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1569] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1570] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1571] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1572] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1573] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1574] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1575] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1576] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1577] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1578] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1579] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1580] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1581] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1582] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1583] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1584] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1585] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1586] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1587] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1588] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1589] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1590] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1591] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1592] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1593] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1594] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1595] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1596] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1597] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1598] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1599] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1600] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1601] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1602] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1603] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1604] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1605] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1606] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1607] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1608] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1609] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1610] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1611] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1612] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1613] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1614] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1615] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1616] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1617] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1618] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1619] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1620] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1621] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1622] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1623] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1624] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1625] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1626] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1627] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1628] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1629] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1630] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1631] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[1632] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1633] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1634] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1635] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1636] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1637] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1638] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1639] = s[0] ? pos_SNs[89] : pos_SNs[89];
	assign level0[1640] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1641] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1642] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1643] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1644] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1645] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1646] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1647] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1648] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1649] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1650] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1651] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1652] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1653] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1654] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1655] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1656] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1657] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1658] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1659] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1660] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1661] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1662] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1663] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1664] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1665] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1666] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1667] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1668] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1669] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1670] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1671] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1672] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1673] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1674] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1675] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1676] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1677] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1678] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1679] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[1680] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1681] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1682] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1683] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1684] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1685] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1686] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1687] = s[0] ? pos_SNs[101] : pos_SNs[101];
	assign level0[1688] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1689] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1690] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1691] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1692] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1693] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1694] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1695] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[1696] = s[0] ? neg_SNs[37] : neg_SNs[37];
	assign level0[1697] = s[0] ? neg_SNs[37] : neg_SNs[37];
	assign level0[1698] = s[0] ? neg_SNs[37] : neg_SNs[37];
	assign level0[1699] = s[0] ? neg_SNs[37] : neg_SNs[37];
	assign level0[1700] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1701] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1702] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1703] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1704] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[1705] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[1706] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[1707] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[1708] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1709] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1710] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1711] = s[0] ? pos_SNs[40] : pos_SNs[40];
	assign level0[1712] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1713] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1714] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1715] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1716] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1717] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1718] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1719] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1720] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1721] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1722] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1723] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1724] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1725] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1726] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1727] = s[0] ? pos_SNs[49] : pos_SNs[49];
	assign level0[1728] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1729] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1730] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1731] = s[0] ? neg_SNs[51] : neg_SNs[51];
	assign level0[1732] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1733] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1734] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1735] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1736] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1737] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1738] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1739] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1740] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1741] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1742] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1743] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1744] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1745] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1746] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1747] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[1748] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1749] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1750] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1751] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1752] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1753] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1754] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1755] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1756] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1757] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1758] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1759] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1760] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1761] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1762] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1763] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1764] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1765] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1766] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1767] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[1768] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1769] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1770] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1771] = s[0] ? pos_SNs[68] : pos_SNs[68];
	assign level0[1772] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1773] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1774] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1775] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1776] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1777] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1778] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1779] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1780] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1781] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1782] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1783] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1784] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1785] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1786] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1787] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1788] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1789] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1790] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1791] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1792] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1793] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1794] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1795] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1796] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1797] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1798] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1799] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1800] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1801] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1802] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1803] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1804] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1805] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1806] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1807] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1808] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1809] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1810] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1811] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[1812] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1813] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1814] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1815] = s[0] ? neg_SNs[81] : neg_SNs[81];
	assign level0[1816] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1817] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1818] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1819] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1820] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1821] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1822] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1823] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1824] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1825] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1826] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1827] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1828] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1829] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1830] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1831] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1832] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1833] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1834] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1835] = s[0] ? pos_SNs[92] : pos_SNs[92];
	assign level0[1836] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1837] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1838] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1839] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1840] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1841] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1842] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1843] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1844] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1845] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1846] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1847] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[1848] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1849] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1850] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1851] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[1852] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1853] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1854] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1855] = s[0] ? pos_SNs[99] : pos_SNs[99];
	assign level0[1856] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1857] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1858] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1859] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1860] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1861] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1862] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1863] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1864] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1865] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1866] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1867] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[1868] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1869] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1870] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1871] = s[0] ? pos_SNs[108] : pos_SNs[108];
	assign level0[1872] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[1873] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[1874] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[1875] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[1876] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1877] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1878] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1879] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[1880] = s[0] ? neg_SNs[111] : neg_SNs[111];
	assign level0[1881] = s[0] ? neg_SNs[111] : neg_SNs[111];
	assign level0[1882] = s[0] ? neg_SNs[111] : neg_SNs[111];
	assign level0[1883] = s[0] ? neg_SNs[111] : neg_SNs[111];
	assign level0[1884] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1885] = s[0] ? pos_SNs[29] : pos_SNs[29];
	assign level0[1886] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1887] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[1888] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1889] = s[0] ? pos_SNs[31] : pos_SNs[31];
	assign level0[1890] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1891] = s[0] ? neg_SNs[32] : neg_SNs[32];
	assign level0[1892] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1893] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1894] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1895] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[1896] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1897] = s[0] ? pos_SNs[43] : pos_SNs[43];
	assign level0[1898] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1899] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1900] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1901] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1902] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1903] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1904] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1905] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1906] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1907] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1908] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1909] = s[0] ? pos_SNs[63] : pos_SNs[63];
	assign level0[1910] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1911] = s[0] ? neg_SNs[64] : neg_SNs[64];
	assign level0[1912] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1913] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1914] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1915] = s[0] ? neg_SNs[69] : neg_SNs[69];
	assign level0[1916] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1917] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1918] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1919] = s[0] ? neg_SNs[71] : neg_SNs[71];
	assign level0[1920] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1921] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1922] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1923] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1924] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1925] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1926] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1927] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1928] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1929] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1930] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1931] = s[0] ? neg_SNs[77] : neg_SNs[77];
	assign level0[1932] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1933] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1934] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1935] = s[0] ? neg_SNs[79] : neg_SNs[79];
	assign level0[1936] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1937] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1938] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1939] = s[0] ? neg_SNs[84] : neg_SNs[84];
	assign level0[1940] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1941] = s[0] ? pos_SNs[85] : pos_SNs[85];
	assign level0[1942] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1943] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1944] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1945] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[1946] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1947] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[1948] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1949] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[1950] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1951] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[1952] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1953] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[1954] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1955] = s[0] ? neg_SNs[107] : neg_SNs[107];
	assign level0[1956] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1957] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[1958] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1959] = s[0] ? neg_SNs[116] : neg_SNs[116];
	assign level0[1960] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1961] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[1962] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1963] = s[0] ? neg_SNs[118] : neg_SNs[118];
	assign level0[1964] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1965] = s[0] ? pos_SNs[119] : pos_SNs[119];
	assign level0[1966] = s[0] ? neg_SNs[21] : neg_SNs[21];
	assign level0[1967] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[1968] = s[0] ? neg_SNs[23] : neg_SNs[23];
	assign level0[1969] = s[0] ? pos_SNs[24] : pos_SNs[24];
	assign level0[1970] = s[0] ? pos_SNs[27] : pos_SNs[27];
	assign level0[1971] = s[0] ? neg_SNs[28] : neg_SNs[28];
	assign level0[1972] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[1973] = s[0] ? neg_SNs[35] : neg_SNs[35];
	assign level0[1974] = s[0] ? pos_SNs[36] : pos_SNs[36];
	assign level0[1975] = s[0] ? pos_SNs[38] : pos_SNs[38];
	assign level0[1976] = s[0] ? neg_SNs[39] : neg_SNs[39];
	assign level0[1977] = s[0] ? neg_SNs[44] : neg_SNs[44];
	assign level0[1978] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[1979] = s[0] ? neg_SNs[48] : neg_SNs[48];
	assign level0[1980] = s[0] ? pos_SNs[52] : pos_SNs[52];
	assign level0[1981] = s[0] ? neg_SNs[53] : neg_SNs[53];
	assign level0[1982] = s[0] ? pos_SNs[54] : pos_SNs[54];
	assign level0[1983] = s[0] ? neg_SNs[55] : neg_SNs[55];
	assign level0[1984] = s[0] ? neg_SNs[57] : neg_SNs[57];
	assign level0[1985] = s[0] ? neg_SNs[60] : neg_SNs[60];
	assign level0[1986] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[1987] = s[0] ? pos_SNs[65] : pos_SNs[65];
	assign level0[1988] = s[0] ? pos_SNs[70] : pos_SNs[70];
	assign level0[1989] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[1990] = s[0] ? neg_SNs[73] : neg_SNs[73];
	assign level0[1991] = s[0] ? pos_SNs[74] : pos_SNs[74];
	assign level0[1992] = s[0] ? neg_SNs[75] : neg_SNs[75];
	assign level0[1993] = s[0] ? pos_SNs[76] : pos_SNs[76];
	assign level0[1994] = s[0] ? pos_SNs[78] : pos_SNs[78];
	assign level0[1995] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[1996] = s[0] ? neg_SNs[86] : neg_SNs[86];
	assign level0[1997] = s[0] ? neg_SNs[88] : neg_SNs[88];
	assign level0[1998] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[1999] = s[0] ? neg_SNs[93] : neg_SNs[93];
	assign level0[2000] = s[0] ? pos_SNs[94] : pos_SNs[94];
	assign level0[2001] = s[0] ? neg_SNs[95] : neg_SNs[95];
	assign level0[2002] = s[0] ? pos_SNs[96] : pos_SNs[96];
	assign level0[2003] = s[0] ? neg_SNs[100] : neg_SNs[100];
	assign level0[2004] = s[0] ? pos_SNs[103] : pos_SNs[103];
	assign level0[2005] = s[0] ? neg_SNs[104] : neg_SNs[104];
	assign level0[2006] = s[0] ? neg_SNs[109] : neg_SNs[109];
	assign level0[2007] = s[0] ? pos_SNs[110] : pos_SNs[110];
	assign level0[2008] = s[0] ? pos_SNs[112] : pos_SNs[112];
	assign level0[2009] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[2010] = s[0] ? pos_SNs[115] : pos_SNs[115];
	assign level0[2011] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[2012] = s[0] ? pos_SNs[121] : pos_SNs[121];
	assign level0[2013] = s[0] ? pos_SNs[124] : pos_SNs[124];
	assign level0[2014] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[2015] = s[0] ? pos_SNs[126] : pos_SNs[126];
	assign level0[2016] = s[0] ? neg_SNs[127] : neg_SNs[127];
	assign level0[2017] = s[0] ? neg_SNs[12] : neg_SNs[12];
	assign level0[2018] = s[0] ? neg_SNs[14] : neg_SNs[14];
	assign level0[2019] = s[0] ? neg_SNs[16] : neg_SNs[16];
	assign level0[2020] = s[0] ? neg_SNs[19] : neg_SNs[19];
	assign level0[2021] = s[0] ? pos_SNs[22] : pos_SNs[22];
	assign level0[2022] = s[0] ? neg_SNs[25] : neg_SNs[25];
	assign level0[2023] = s[0] ? neg_SNs[30] : neg_SNs[30];
	assign level0[2024] = s[0] ? pos_SNs[33] : pos_SNs[33];
	assign level0[2025] = s[0] ? neg_SNs[41] : neg_SNs[41];
	assign level0[2026] = s[0] ? pos_SNs[45] : pos_SNs[45];
	assign level0[2027] = s[0] ? pos_SNs[47] : pos_SNs[47];
	assign level0[2028] = s[0] ? pos_SNs[56] : pos_SNs[56];
	assign level0[2029] = s[0] ? pos_SNs[59] : pos_SNs[59];
	assign level0[2030] = s[0] ? neg_SNs[62] : neg_SNs[62];
	assign level0[2031] = s[0] ? neg_SNs[67] : neg_SNs[67];
	assign level0[2032] = s[0] ? pos_SNs[72] : pos_SNs[72];
	assign level0[2033] = s[0] ? pos_SNs[80] : pos_SNs[80];
	assign level0[2034] = s[0] ? pos_SNs[83] : pos_SNs[83];
	assign level0[2035] = s[0] ? pos_SNs[87] : pos_SNs[87];
	assign level0[2036] = s[0] ? neg_SNs[91] : neg_SNs[91];
	assign level0[2037] = s[0] ? neg_SNs[97] : neg_SNs[97];
	assign level0[2038] = s[0] ? neg_SNs[102] : neg_SNs[102];
	assign level0[2039] = s[0] ? pos_SNs[105] : pos_SNs[105];
	assign level0[2040] = s[0] ? neg_SNs[113] : neg_SNs[113];
	assign level0[2041] = s[0] ? pos_SNs[117] : pos_SNs[117];
	assign level0[2042] = s[0] ? neg_SNs[120] : neg_SNs[120];
	assign level0[2043] = s[0] ? neg_SNs[125] : neg_SNs[125];
	assign level0[2044] = s[0] ? pos_SNs[128] : pos_SNs[128];
	assign level0[2045] = s[0] ? pos_SNs[131] : pos_SNs[131];
	assign level0[2046] = s[0] ? pos_SNs[133] : pos_SNs[133];
	assign level0[2047] = s[0] ? pos_SNs[135] : pos_SNs[135];

	assign level1[0] = s[1] ? level0[0] : level0[1];
	assign level1[1] = s[1] ? level0[2] : level0[3];
	assign level1[2] = s[1] ? level0[4] : level0[5];
	assign level1[3] = s[1] ? level0[6] : level0[7];
	assign level1[4] = s[1] ? level0[8] : level0[9];
	assign level1[5] = s[1] ? level0[10] : level0[11];
	assign level1[6] = s[1] ? level0[12] : level0[13];
	assign level1[7] = s[1] ? level0[14] : level0[15];
	assign level1[8] = s[1] ? level0[16] : level0[17];
	assign level1[9] = s[1] ? level0[18] : level0[19];
	assign level1[10] = s[1] ? level0[20] : level0[21];
	assign level1[11] = s[1] ? level0[22] : level0[23];
	assign level1[12] = s[1] ? level0[24] : level0[25];
	assign level1[13] = s[1] ? level0[26] : level0[27];
	assign level1[14] = s[1] ? level0[28] : level0[29];
	assign level1[15] = s[1] ? level0[30] : level0[31];
	assign level1[16] = s[1] ? level0[32] : level0[33];
	assign level1[17] = s[1] ? level0[34] : level0[35];
	assign level1[18] = s[1] ? level0[36] : level0[37];
	assign level1[19] = s[1] ? level0[38] : level0[39];
	assign level1[20] = s[1] ? level0[40] : level0[41];
	assign level1[21] = s[1] ? level0[42] : level0[43];
	assign level1[22] = s[1] ? level0[44] : level0[45];
	assign level1[23] = s[1] ? level0[46] : level0[47];
	assign level1[24] = s[1] ? level0[48] : level0[49];
	assign level1[25] = s[1] ? level0[50] : level0[51];
	assign level1[26] = s[1] ? level0[52] : level0[53];
	assign level1[27] = s[1] ? level0[54] : level0[55];
	assign level1[28] = s[1] ? level0[56] : level0[57];
	assign level1[29] = s[1] ? level0[58] : level0[59];
	assign level1[30] = s[1] ? level0[60] : level0[61];
	assign level1[31] = s[1] ? level0[62] : level0[63];
	assign level1[32] = s[1] ? level0[64] : level0[65];
	assign level1[33] = s[1] ? level0[66] : level0[67];
	assign level1[34] = s[1] ? level0[68] : level0[69];
	assign level1[35] = s[1] ? level0[70] : level0[71];
	assign level1[36] = s[1] ? level0[72] : level0[73];
	assign level1[37] = s[1] ? level0[74] : level0[75];
	assign level1[38] = s[1] ? level0[76] : level0[77];
	assign level1[39] = s[1] ? level0[78] : level0[79];
	assign level1[40] = s[1] ? level0[80] : level0[81];
	assign level1[41] = s[1] ? level0[82] : level0[83];
	assign level1[42] = s[1] ? level0[84] : level0[85];
	assign level1[43] = s[1] ? level0[86] : level0[87];
	assign level1[44] = s[1] ? level0[88] : level0[89];
	assign level1[45] = s[1] ? level0[90] : level0[91];
	assign level1[46] = s[1] ? level0[92] : level0[93];
	assign level1[47] = s[1] ? level0[94] : level0[95];
	assign level1[48] = s[1] ? level0[96] : level0[97];
	assign level1[49] = s[1] ? level0[98] : level0[99];
	assign level1[50] = s[1] ? level0[100] : level0[101];
	assign level1[51] = s[1] ? level0[102] : level0[103];
	assign level1[52] = s[1] ? level0[104] : level0[105];
	assign level1[53] = s[1] ? level0[106] : level0[107];
	assign level1[54] = s[1] ? level0[108] : level0[109];
	assign level1[55] = s[1] ? level0[110] : level0[111];
	assign level1[56] = s[1] ? level0[112] : level0[113];
	assign level1[57] = s[1] ? level0[114] : level0[115];
	assign level1[58] = s[1] ? level0[116] : level0[117];
	assign level1[59] = s[1] ? level0[118] : level0[119];
	assign level1[60] = s[1] ? level0[120] : level0[121];
	assign level1[61] = s[1] ? level0[122] : level0[123];
	assign level1[62] = s[1] ? level0[124] : level0[125];
	assign level1[63] = s[1] ? level0[126] : level0[127];
	assign level1[64] = s[1] ? level0[128] : level0[129];
	assign level1[65] = s[1] ? level0[130] : level0[131];
	assign level1[66] = s[1] ? level0[132] : level0[133];
	assign level1[67] = s[1] ? level0[134] : level0[135];
	assign level1[68] = s[1] ? level0[136] : level0[137];
	assign level1[69] = s[1] ? level0[138] : level0[139];
	assign level1[70] = s[1] ? level0[140] : level0[141];
	assign level1[71] = s[1] ? level0[142] : level0[143];
	assign level1[72] = s[1] ? level0[144] : level0[145];
	assign level1[73] = s[1] ? level0[146] : level0[147];
	assign level1[74] = s[1] ? level0[148] : level0[149];
	assign level1[75] = s[1] ? level0[150] : level0[151];
	assign level1[76] = s[1] ? level0[152] : level0[153];
	assign level1[77] = s[1] ? level0[154] : level0[155];
	assign level1[78] = s[1] ? level0[156] : level0[157];
	assign level1[79] = s[1] ? level0[158] : level0[159];
	assign level1[80] = s[1] ? level0[160] : level0[161];
	assign level1[81] = s[1] ? level0[162] : level0[163];
	assign level1[82] = s[1] ? level0[164] : level0[165];
	assign level1[83] = s[1] ? level0[166] : level0[167];
	assign level1[84] = s[1] ? level0[168] : level0[169];
	assign level1[85] = s[1] ? level0[170] : level0[171];
	assign level1[86] = s[1] ? level0[172] : level0[173];
	assign level1[87] = s[1] ? level0[174] : level0[175];
	assign level1[88] = s[1] ? level0[176] : level0[177];
	assign level1[89] = s[1] ? level0[178] : level0[179];
	assign level1[90] = s[1] ? level0[180] : level0[181];
	assign level1[91] = s[1] ? level0[182] : level0[183];
	assign level1[92] = s[1] ? level0[184] : level0[185];
	assign level1[93] = s[1] ? level0[186] : level0[187];
	assign level1[94] = s[1] ? level0[188] : level0[189];
	assign level1[95] = s[1] ? level0[190] : level0[191];
	assign level1[96] = s[1] ? level0[192] : level0[193];
	assign level1[97] = s[1] ? level0[194] : level0[195];
	assign level1[98] = s[1] ? level0[196] : level0[197];
	assign level1[99] = s[1] ? level0[198] : level0[199];
	assign level1[100] = s[1] ? level0[200] : level0[201];
	assign level1[101] = s[1] ? level0[202] : level0[203];
	assign level1[102] = s[1] ? level0[204] : level0[205];
	assign level1[103] = s[1] ? level0[206] : level0[207];
	assign level1[104] = s[1] ? level0[208] : level0[209];
	assign level1[105] = s[1] ? level0[210] : level0[211];
	assign level1[106] = s[1] ? level0[212] : level0[213];
	assign level1[107] = s[1] ? level0[214] : level0[215];
	assign level1[108] = s[1] ? level0[216] : level0[217];
	assign level1[109] = s[1] ? level0[218] : level0[219];
	assign level1[110] = s[1] ? level0[220] : level0[221];
	assign level1[111] = s[1] ? level0[222] : level0[223];
	assign level1[112] = s[1] ? level0[224] : level0[225];
	assign level1[113] = s[1] ? level0[226] : level0[227];
	assign level1[114] = s[1] ? level0[228] : level0[229];
	assign level1[115] = s[1] ? level0[230] : level0[231];
	assign level1[116] = s[1] ? level0[232] : level0[233];
	assign level1[117] = s[1] ? level0[234] : level0[235];
	assign level1[118] = s[1] ? level0[236] : level0[237];
	assign level1[119] = s[1] ? level0[238] : level0[239];
	assign level1[120] = s[1] ? level0[240] : level0[241];
	assign level1[121] = s[1] ? level0[242] : level0[243];
	assign level1[122] = s[1] ? level0[244] : level0[245];
	assign level1[123] = s[1] ? level0[246] : level0[247];
	assign level1[124] = s[1] ? level0[248] : level0[249];
	assign level1[125] = s[1] ? level0[250] : level0[251];
	assign level1[126] = s[1] ? level0[252] : level0[253];
	assign level1[127] = s[1] ? level0[254] : level0[255];
	assign level1[128] = s[1] ? level0[256] : level0[257];
	assign level1[129] = s[1] ? level0[258] : level0[259];
	assign level1[130] = s[1] ? level0[260] : level0[261];
	assign level1[131] = s[1] ? level0[262] : level0[263];
	assign level1[132] = s[1] ? level0[264] : level0[265];
	assign level1[133] = s[1] ? level0[266] : level0[267];
	assign level1[134] = s[1] ? level0[268] : level0[269];
	assign level1[135] = s[1] ? level0[270] : level0[271];
	assign level1[136] = s[1] ? level0[272] : level0[273];
	assign level1[137] = s[1] ? level0[274] : level0[275];
	assign level1[138] = s[1] ? level0[276] : level0[277];
	assign level1[139] = s[1] ? level0[278] : level0[279];
	assign level1[140] = s[1] ? level0[280] : level0[281];
	assign level1[141] = s[1] ? level0[282] : level0[283];
	assign level1[142] = s[1] ? level0[284] : level0[285];
	assign level1[143] = s[1] ? level0[286] : level0[287];
	assign level1[144] = s[1] ? level0[288] : level0[289];
	assign level1[145] = s[1] ? level0[290] : level0[291];
	assign level1[146] = s[1] ? level0[292] : level0[293];
	assign level1[147] = s[1] ? level0[294] : level0[295];
	assign level1[148] = s[1] ? level0[296] : level0[297];
	assign level1[149] = s[1] ? level0[298] : level0[299];
	assign level1[150] = s[1] ? level0[300] : level0[301];
	assign level1[151] = s[1] ? level0[302] : level0[303];
	assign level1[152] = s[1] ? level0[304] : level0[305];
	assign level1[153] = s[1] ? level0[306] : level0[307];
	assign level1[154] = s[1] ? level0[308] : level0[309];
	assign level1[155] = s[1] ? level0[310] : level0[311];
	assign level1[156] = s[1] ? level0[312] : level0[313];
	assign level1[157] = s[1] ? level0[314] : level0[315];
	assign level1[158] = s[1] ? level0[316] : level0[317];
	assign level1[159] = s[1] ? level0[318] : level0[319];
	assign level1[160] = s[1] ? level0[320] : level0[321];
	assign level1[161] = s[1] ? level0[322] : level0[323];
	assign level1[162] = s[1] ? level0[324] : level0[325];
	assign level1[163] = s[1] ? level0[326] : level0[327];
	assign level1[164] = s[1] ? level0[328] : level0[329];
	assign level1[165] = s[1] ? level0[330] : level0[331];
	assign level1[166] = s[1] ? level0[332] : level0[333];
	assign level1[167] = s[1] ? level0[334] : level0[335];
	assign level1[168] = s[1] ? level0[336] : level0[337];
	assign level1[169] = s[1] ? level0[338] : level0[339];
	assign level1[170] = s[1] ? level0[340] : level0[341];
	assign level1[171] = s[1] ? level0[342] : level0[343];
	assign level1[172] = s[1] ? level0[344] : level0[345];
	assign level1[173] = s[1] ? level0[346] : level0[347];
	assign level1[174] = s[1] ? level0[348] : level0[349];
	assign level1[175] = s[1] ? level0[350] : level0[351];
	assign level1[176] = s[1] ? level0[352] : level0[353];
	assign level1[177] = s[1] ? level0[354] : level0[355];
	assign level1[178] = s[1] ? level0[356] : level0[357];
	assign level1[179] = s[1] ? level0[358] : level0[359];
	assign level1[180] = s[1] ? level0[360] : level0[361];
	assign level1[181] = s[1] ? level0[362] : level0[363];
	assign level1[182] = s[1] ? level0[364] : level0[365];
	assign level1[183] = s[1] ? level0[366] : level0[367];
	assign level1[184] = s[1] ? level0[368] : level0[369];
	assign level1[185] = s[1] ? level0[370] : level0[371];
	assign level1[186] = s[1] ? level0[372] : level0[373];
	assign level1[187] = s[1] ? level0[374] : level0[375];
	assign level1[188] = s[1] ? level0[376] : level0[377];
	assign level1[189] = s[1] ? level0[378] : level0[379];
	assign level1[190] = s[1] ? level0[380] : level0[381];
	assign level1[191] = s[1] ? level0[382] : level0[383];
	assign level1[192] = s[1] ? level0[384] : level0[385];
	assign level1[193] = s[1] ? level0[386] : level0[387];
	assign level1[194] = s[1] ? level0[388] : level0[389];
	assign level1[195] = s[1] ? level0[390] : level0[391];
	assign level1[196] = s[1] ? level0[392] : level0[393];
	assign level1[197] = s[1] ? level0[394] : level0[395];
	assign level1[198] = s[1] ? level0[396] : level0[397];
	assign level1[199] = s[1] ? level0[398] : level0[399];
	assign level1[200] = s[1] ? level0[400] : level0[401];
	assign level1[201] = s[1] ? level0[402] : level0[403];
	assign level1[202] = s[1] ? level0[404] : level0[405];
	assign level1[203] = s[1] ? level0[406] : level0[407];
	assign level1[204] = s[1] ? level0[408] : level0[409];
	assign level1[205] = s[1] ? level0[410] : level0[411];
	assign level1[206] = s[1] ? level0[412] : level0[413];
	assign level1[207] = s[1] ? level0[414] : level0[415];
	assign level1[208] = s[1] ? level0[416] : level0[417];
	assign level1[209] = s[1] ? level0[418] : level0[419];
	assign level1[210] = s[1] ? level0[420] : level0[421];
	assign level1[211] = s[1] ? level0[422] : level0[423];
	assign level1[212] = s[1] ? level0[424] : level0[425];
	assign level1[213] = s[1] ? level0[426] : level0[427];
	assign level1[214] = s[1] ? level0[428] : level0[429];
	assign level1[215] = s[1] ? level0[430] : level0[431];
	assign level1[216] = s[1] ? level0[432] : level0[433];
	assign level1[217] = s[1] ? level0[434] : level0[435];
	assign level1[218] = s[1] ? level0[436] : level0[437];
	assign level1[219] = s[1] ? level0[438] : level0[439];
	assign level1[220] = s[1] ? level0[440] : level0[441];
	assign level1[221] = s[1] ? level0[442] : level0[443];
	assign level1[222] = s[1] ? level0[444] : level0[445];
	assign level1[223] = s[1] ? level0[446] : level0[447];
	assign level1[224] = s[1] ? level0[448] : level0[449];
	assign level1[225] = s[1] ? level0[450] : level0[451];
	assign level1[226] = s[1] ? level0[452] : level0[453];
	assign level1[227] = s[1] ? level0[454] : level0[455];
	assign level1[228] = s[1] ? level0[456] : level0[457];
	assign level1[229] = s[1] ? level0[458] : level0[459];
	assign level1[230] = s[1] ? level0[460] : level0[461];
	assign level1[231] = s[1] ? level0[462] : level0[463];
	assign level1[232] = s[1] ? level0[464] : level0[465];
	assign level1[233] = s[1] ? level0[466] : level0[467];
	assign level1[234] = s[1] ? level0[468] : level0[469];
	assign level1[235] = s[1] ? level0[470] : level0[471];
	assign level1[236] = s[1] ? level0[472] : level0[473];
	assign level1[237] = s[1] ? level0[474] : level0[475];
	assign level1[238] = s[1] ? level0[476] : level0[477];
	assign level1[239] = s[1] ? level0[478] : level0[479];
	assign level1[240] = s[1] ? level0[480] : level0[481];
	assign level1[241] = s[1] ? level0[482] : level0[483];
	assign level1[242] = s[1] ? level0[484] : level0[485];
	assign level1[243] = s[1] ? level0[486] : level0[487];
	assign level1[244] = s[1] ? level0[488] : level0[489];
	assign level1[245] = s[1] ? level0[490] : level0[491];
	assign level1[246] = s[1] ? level0[492] : level0[493];
	assign level1[247] = s[1] ? level0[494] : level0[495];
	assign level1[248] = s[1] ? level0[496] : level0[497];
	assign level1[249] = s[1] ? level0[498] : level0[499];
	assign level1[250] = s[1] ? level0[500] : level0[501];
	assign level1[251] = s[1] ? level0[502] : level0[503];
	assign level1[252] = s[1] ? level0[504] : level0[505];
	assign level1[253] = s[1] ? level0[506] : level0[507];
	assign level1[254] = s[1] ? level0[508] : level0[509];
	assign level1[255] = s[1] ? level0[510] : level0[511];
	assign level1[256] = s[1] ? level0[512] : level0[513];
	assign level1[257] = s[1] ? level0[514] : level0[515];
	assign level1[258] = s[1] ? level0[516] : level0[517];
	assign level1[259] = s[1] ? level0[518] : level0[519];
	assign level1[260] = s[1] ? level0[520] : level0[521];
	assign level1[261] = s[1] ? level0[522] : level0[523];
	assign level1[262] = s[1] ? level0[524] : level0[525];
	assign level1[263] = s[1] ? level0[526] : level0[527];
	assign level1[264] = s[1] ? level0[528] : level0[529];
	assign level1[265] = s[1] ? level0[530] : level0[531];
	assign level1[266] = s[1] ? level0[532] : level0[533];
	assign level1[267] = s[1] ? level0[534] : level0[535];
	assign level1[268] = s[1] ? level0[536] : level0[537];
	assign level1[269] = s[1] ? level0[538] : level0[539];
	assign level1[270] = s[1] ? level0[540] : level0[541];
	assign level1[271] = s[1] ? level0[542] : level0[543];
	assign level1[272] = s[1] ? level0[544] : level0[545];
	assign level1[273] = s[1] ? level0[546] : level0[547];
	assign level1[274] = s[1] ? level0[548] : level0[549];
	assign level1[275] = s[1] ? level0[550] : level0[551];
	assign level1[276] = s[1] ? level0[552] : level0[553];
	assign level1[277] = s[1] ? level0[554] : level0[555];
	assign level1[278] = s[1] ? level0[556] : level0[557];
	assign level1[279] = s[1] ? level0[558] : level0[559];
	assign level1[280] = s[1] ? level0[560] : level0[561];
	assign level1[281] = s[1] ? level0[562] : level0[563];
	assign level1[282] = s[1] ? level0[564] : level0[565];
	assign level1[283] = s[1] ? level0[566] : level0[567];
	assign level1[284] = s[1] ? level0[568] : level0[569];
	assign level1[285] = s[1] ? level0[570] : level0[571];
	assign level1[286] = s[1] ? level0[572] : level0[573];
	assign level1[287] = s[1] ? level0[574] : level0[575];
	assign level1[288] = s[1] ? level0[576] : level0[577];
	assign level1[289] = s[1] ? level0[578] : level0[579];
	assign level1[290] = s[1] ? level0[580] : level0[581];
	assign level1[291] = s[1] ? level0[582] : level0[583];
	assign level1[292] = s[1] ? level0[584] : level0[585];
	assign level1[293] = s[1] ? level0[586] : level0[587];
	assign level1[294] = s[1] ? level0[588] : level0[589];
	assign level1[295] = s[1] ? level0[590] : level0[591];
	assign level1[296] = s[1] ? level0[592] : level0[593];
	assign level1[297] = s[1] ? level0[594] : level0[595];
	assign level1[298] = s[1] ? level0[596] : level0[597];
	assign level1[299] = s[1] ? level0[598] : level0[599];
	assign level1[300] = s[1] ? level0[600] : level0[601];
	assign level1[301] = s[1] ? level0[602] : level0[603];
	assign level1[302] = s[1] ? level0[604] : level0[605];
	assign level1[303] = s[1] ? level0[606] : level0[607];
	assign level1[304] = s[1] ? level0[608] : level0[609];
	assign level1[305] = s[1] ? level0[610] : level0[611];
	assign level1[306] = s[1] ? level0[612] : level0[613];
	assign level1[307] = s[1] ? level0[614] : level0[615];
	assign level1[308] = s[1] ? level0[616] : level0[617];
	assign level1[309] = s[1] ? level0[618] : level0[619];
	assign level1[310] = s[1] ? level0[620] : level0[621];
	assign level1[311] = s[1] ? level0[622] : level0[623];
	assign level1[312] = s[1] ? level0[624] : level0[625];
	assign level1[313] = s[1] ? level0[626] : level0[627];
	assign level1[314] = s[1] ? level0[628] : level0[629];
	assign level1[315] = s[1] ? level0[630] : level0[631];
	assign level1[316] = s[1] ? level0[632] : level0[633];
	assign level1[317] = s[1] ? level0[634] : level0[635];
	assign level1[318] = s[1] ? level0[636] : level0[637];
	assign level1[319] = s[1] ? level0[638] : level0[639];
	assign level1[320] = s[1] ? level0[640] : level0[641];
	assign level1[321] = s[1] ? level0[642] : level0[643];
	assign level1[322] = s[1] ? level0[644] : level0[645];
	assign level1[323] = s[1] ? level0[646] : level0[647];
	assign level1[324] = s[1] ? level0[648] : level0[649];
	assign level1[325] = s[1] ? level0[650] : level0[651];
	assign level1[326] = s[1] ? level0[652] : level0[653];
	assign level1[327] = s[1] ? level0[654] : level0[655];
	assign level1[328] = s[1] ? level0[656] : level0[657];
	assign level1[329] = s[1] ? level0[658] : level0[659];
	assign level1[330] = s[1] ? level0[660] : level0[661];
	assign level1[331] = s[1] ? level0[662] : level0[663];
	assign level1[332] = s[1] ? level0[664] : level0[665];
	assign level1[333] = s[1] ? level0[666] : level0[667];
	assign level1[334] = s[1] ? level0[668] : level0[669];
	assign level1[335] = s[1] ? level0[670] : level0[671];
	assign level1[336] = s[1] ? level0[672] : level0[673];
	assign level1[337] = s[1] ? level0[674] : level0[675];
	assign level1[338] = s[1] ? level0[676] : level0[677];
	assign level1[339] = s[1] ? level0[678] : level0[679];
	assign level1[340] = s[1] ? level0[680] : level0[681];
	assign level1[341] = s[1] ? level0[682] : level0[683];
	assign level1[342] = s[1] ? level0[684] : level0[685];
	assign level1[343] = s[1] ? level0[686] : level0[687];
	assign level1[344] = s[1] ? level0[688] : level0[689];
	assign level1[345] = s[1] ? level0[690] : level0[691];
	assign level1[346] = s[1] ? level0[692] : level0[693];
	assign level1[347] = s[1] ? level0[694] : level0[695];
	assign level1[348] = s[1] ? level0[696] : level0[697];
	assign level1[349] = s[1] ? level0[698] : level0[699];
	assign level1[350] = s[1] ? level0[700] : level0[701];
	assign level1[351] = s[1] ? level0[702] : level0[703];
	assign level1[352] = s[1] ? level0[704] : level0[705];
	assign level1[353] = s[1] ? level0[706] : level0[707];
	assign level1[354] = s[1] ? level0[708] : level0[709];
	assign level1[355] = s[1] ? level0[710] : level0[711];
	assign level1[356] = s[1] ? level0[712] : level0[713];
	assign level1[357] = s[1] ? level0[714] : level0[715];
	assign level1[358] = s[1] ? level0[716] : level0[717];
	assign level1[359] = s[1] ? level0[718] : level0[719];
	assign level1[360] = s[1] ? level0[720] : level0[721];
	assign level1[361] = s[1] ? level0[722] : level0[723];
	assign level1[362] = s[1] ? level0[724] : level0[725];
	assign level1[363] = s[1] ? level0[726] : level0[727];
	assign level1[364] = s[1] ? level0[728] : level0[729];
	assign level1[365] = s[1] ? level0[730] : level0[731];
	assign level1[366] = s[1] ? level0[732] : level0[733];
	assign level1[367] = s[1] ? level0[734] : level0[735];
	assign level1[368] = s[1] ? level0[736] : level0[737];
	assign level1[369] = s[1] ? level0[738] : level0[739];
	assign level1[370] = s[1] ? level0[740] : level0[741];
	assign level1[371] = s[1] ? level0[742] : level0[743];
	assign level1[372] = s[1] ? level0[744] : level0[745];
	assign level1[373] = s[1] ? level0[746] : level0[747];
	assign level1[374] = s[1] ? level0[748] : level0[749];
	assign level1[375] = s[1] ? level0[750] : level0[751];
	assign level1[376] = s[1] ? level0[752] : level0[753];
	assign level1[377] = s[1] ? level0[754] : level0[755];
	assign level1[378] = s[1] ? level0[756] : level0[757];
	assign level1[379] = s[1] ? level0[758] : level0[759];
	assign level1[380] = s[1] ? level0[760] : level0[761];
	assign level1[381] = s[1] ? level0[762] : level0[763];
	assign level1[382] = s[1] ? level0[764] : level0[765];
	assign level1[383] = s[1] ? level0[766] : level0[767];
	assign level1[384] = s[1] ? level0[768] : level0[769];
	assign level1[385] = s[1] ? level0[770] : level0[771];
	assign level1[386] = s[1] ? level0[772] : level0[773];
	assign level1[387] = s[1] ? level0[774] : level0[775];
	assign level1[388] = s[1] ? level0[776] : level0[777];
	assign level1[389] = s[1] ? level0[778] : level0[779];
	assign level1[390] = s[1] ? level0[780] : level0[781];
	assign level1[391] = s[1] ? level0[782] : level0[783];
	assign level1[392] = s[1] ? level0[784] : level0[785];
	assign level1[393] = s[1] ? level0[786] : level0[787];
	assign level1[394] = s[1] ? level0[788] : level0[789];
	assign level1[395] = s[1] ? level0[790] : level0[791];
	assign level1[396] = s[1] ? level0[792] : level0[793];
	assign level1[397] = s[1] ? level0[794] : level0[795];
	assign level1[398] = s[1] ? level0[796] : level0[797];
	assign level1[399] = s[1] ? level0[798] : level0[799];
	assign level1[400] = s[1] ? level0[800] : level0[801];
	assign level1[401] = s[1] ? level0[802] : level0[803];
	assign level1[402] = s[1] ? level0[804] : level0[805];
	assign level1[403] = s[1] ? level0[806] : level0[807];
	assign level1[404] = s[1] ? level0[808] : level0[809];
	assign level1[405] = s[1] ? level0[810] : level0[811];
	assign level1[406] = s[1] ? level0[812] : level0[813];
	assign level1[407] = s[1] ? level0[814] : level0[815];
	assign level1[408] = s[1] ? level0[816] : level0[817];
	assign level1[409] = s[1] ? level0[818] : level0[819];
	assign level1[410] = s[1] ? level0[820] : level0[821];
	assign level1[411] = s[1] ? level0[822] : level0[823];
	assign level1[412] = s[1] ? level0[824] : level0[825];
	assign level1[413] = s[1] ? level0[826] : level0[827];
	assign level1[414] = s[1] ? level0[828] : level0[829];
	assign level1[415] = s[1] ? level0[830] : level0[831];
	assign level1[416] = s[1] ? level0[832] : level0[833];
	assign level1[417] = s[1] ? level0[834] : level0[835];
	assign level1[418] = s[1] ? level0[836] : level0[837];
	assign level1[419] = s[1] ? level0[838] : level0[839];
	assign level1[420] = s[1] ? level0[840] : level0[841];
	assign level1[421] = s[1] ? level0[842] : level0[843];
	assign level1[422] = s[1] ? level0[844] : level0[845];
	assign level1[423] = s[1] ? level0[846] : level0[847];
	assign level1[424] = s[1] ? level0[848] : level0[849];
	assign level1[425] = s[1] ? level0[850] : level0[851];
	assign level1[426] = s[1] ? level0[852] : level0[853];
	assign level1[427] = s[1] ? level0[854] : level0[855];
	assign level1[428] = s[1] ? level0[856] : level0[857];
	assign level1[429] = s[1] ? level0[858] : level0[859];
	assign level1[430] = s[1] ? level0[860] : level0[861];
	assign level1[431] = s[1] ? level0[862] : level0[863];
	assign level1[432] = s[1] ? level0[864] : level0[865];
	assign level1[433] = s[1] ? level0[866] : level0[867];
	assign level1[434] = s[1] ? level0[868] : level0[869];
	assign level1[435] = s[1] ? level0[870] : level0[871];
	assign level1[436] = s[1] ? level0[872] : level0[873];
	assign level1[437] = s[1] ? level0[874] : level0[875];
	assign level1[438] = s[1] ? level0[876] : level0[877];
	assign level1[439] = s[1] ? level0[878] : level0[879];
	assign level1[440] = s[1] ? level0[880] : level0[881];
	assign level1[441] = s[1] ? level0[882] : level0[883];
	assign level1[442] = s[1] ? level0[884] : level0[885];
	assign level1[443] = s[1] ? level0[886] : level0[887];
	assign level1[444] = s[1] ? level0[888] : level0[889];
	assign level1[445] = s[1] ? level0[890] : level0[891];
	assign level1[446] = s[1] ? level0[892] : level0[893];
	assign level1[447] = s[1] ? level0[894] : level0[895];
	assign level1[448] = s[1] ? level0[896] : level0[897];
	assign level1[449] = s[1] ? level0[898] : level0[899];
	assign level1[450] = s[1] ? level0[900] : level0[901];
	assign level1[451] = s[1] ? level0[902] : level0[903];
	assign level1[452] = s[1] ? level0[904] : level0[905];
	assign level1[453] = s[1] ? level0[906] : level0[907];
	assign level1[454] = s[1] ? level0[908] : level0[909];
	assign level1[455] = s[1] ? level0[910] : level0[911];
	assign level1[456] = s[1] ? level0[912] : level0[913];
	assign level1[457] = s[1] ? level0[914] : level0[915];
	assign level1[458] = s[1] ? level0[916] : level0[917];
	assign level1[459] = s[1] ? level0[918] : level0[919];
	assign level1[460] = s[1] ? level0[920] : level0[921];
	assign level1[461] = s[1] ? level0[922] : level0[923];
	assign level1[462] = s[1] ? level0[924] : level0[925];
	assign level1[463] = s[1] ? level0[926] : level0[927];
	assign level1[464] = s[1] ? level0[928] : level0[929];
	assign level1[465] = s[1] ? level0[930] : level0[931];
	assign level1[466] = s[1] ? level0[932] : level0[933];
	assign level1[467] = s[1] ? level0[934] : level0[935];
	assign level1[468] = s[1] ? level0[936] : level0[937];
	assign level1[469] = s[1] ? level0[938] : level0[939];
	assign level1[470] = s[1] ? level0[940] : level0[941];
	assign level1[471] = s[1] ? level0[942] : level0[943];
	assign level1[472] = s[1] ? level0[944] : level0[945];
	assign level1[473] = s[1] ? level0[946] : level0[947];
	assign level1[474] = s[1] ? level0[948] : level0[949];
	assign level1[475] = s[1] ? level0[950] : level0[951];
	assign level1[476] = s[1] ? level0[952] : level0[953];
	assign level1[477] = s[1] ? level0[954] : level0[955];
	assign level1[478] = s[1] ? level0[956] : level0[957];
	assign level1[479] = s[1] ? level0[958] : level0[959];
	assign level1[480] = s[1] ? level0[960] : level0[961];
	assign level1[481] = s[1] ? level0[962] : level0[963];
	assign level1[482] = s[1] ? level0[964] : level0[965];
	assign level1[483] = s[1] ? level0[966] : level0[967];
	assign level1[484] = s[1] ? level0[968] : level0[969];
	assign level1[485] = s[1] ? level0[970] : level0[971];
	assign level1[486] = s[1] ? level0[972] : level0[973];
	assign level1[487] = s[1] ? level0[974] : level0[975];
	assign level1[488] = s[1] ? level0[976] : level0[977];
	assign level1[489] = s[1] ? level0[978] : level0[979];
	assign level1[490] = s[1] ? level0[980] : level0[981];
	assign level1[491] = s[1] ? level0[982] : level0[983];
	assign level1[492] = s[1] ? level0[984] : level0[985];
	assign level1[493] = s[1] ? level0[986] : level0[987];
	assign level1[494] = s[1] ? level0[988] : level0[989];
	assign level1[495] = s[1] ? level0[990] : level0[991];
	assign level1[496] = s[1] ? level0[992] : level0[993];
	assign level1[497] = s[1] ? level0[994] : level0[995];
	assign level1[498] = s[1] ? level0[996] : level0[997];
	assign level1[499] = s[1] ? level0[998] : level0[999];
	assign level1[500] = s[1] ? level0[1000] : level0[1001];
	assign level1[501] = s[1] ? level0[1002] : level0[1003];
	assign level1[502] = s[1] ? level0[1004] : level0[1005];
	assign level1[503] = s[1] ? level0[1006] : level0[1007];
	assign level1[504] = s[1] ? level0[1008] : level0[1009];
	assign level1[505] = s[1] ? level0[1010] : level0[1011];
	assign level1[506] = s[1] ? level0[1012] : level0[1013];
	assign level1[507] = s[1] ? level0[1014] : level0[1015];
	assign level1[508] = s[1] ? level0[1016] : level0[1017];
	assign level1[509] = s[1] ? level0[1018] : level0[1019];
	assign level1[510] = s[1] ? level0[1020] : level0[1021];
	assign level1[511] = s[1] ? level0[1022] : level0[1023];
	assign level1[512] = s[1] ? level0[1024] : level0[1025];
	assign level1[513] = s[1] ? level0[1026] : level0[1027];
	assign level1[514] = s[1] ? level0[1028] : level0[1029];
	assign level1[515] = s[1] ? level0[1030] : level0[1031];
	assign level1[516] = s[1] ? level0[1032] : level0[1033];
	assign level1[517] = s[1] ? level0[1034] : level0[1035];
	assign level1[518] = s[1] ? level0[1036] : level0[1037];
	assign level1[519] = s[1] ? level0[1038] : level0[1039];
	assign level1[520] = s[1] ? level0[1040] : level0[1041];
	assign level1[521] = s[1] ? level0[1042] : level0[1043];
	assign level1[522] = s[1] ? level0[1044] : level0[1045];
	assign level1[523] = s[1] ? level0[1046] : level0[1047];
	assign level1[524] = s[1] ? level0[1048] : level0[1049];
	assign level1[525] = s[1] ? level0[1050] : level0[1051];
	assign level1[526] = s[1] ? level0[1052] : level0[1053];
	assign level1[527] = s[1] ? level0[1054] : level0[1055];
	assign level1[528] = s[1] ? level0[1056] : level0[1057];
	assign level1[529] = s[1] ? level0[1058] : level0[1059];
	assign level1[530] = s[1] ? level0[1060] : level0[1061];
	assign level1[531] = s[1] ? level0[1062] : level0[1063];
	assign level1[532] = s[1] ? level0[1064] : level0[1065];
	assign level1[533] = s[1] ? level0[1066] : level0[1067];
	assign level1[534] = s[1] ? level0[1068] : level0[1069];
	assign level1[535] = s[1] ? level0[1070] : level0[1071];
	assign level1[536] = s[1] ? level0[1072] : level0[1073];
	assign level1[537] = s[1] ? level0[1074] : level0[1075];
	assign level1[538] = s[1] ? level0[1076] : level0[1077];
	assign level1[539] = s[1] ? level0[1078] : level0[1079];
	assign level1[540] = s[1] ? level0[1080] : level0[1081];
	assign level1[541] = s[1] ? level0[1082] : level0[1083];
	assign level1[542] = s[1] ? level0[1084] : level0[1085];
	assign level1[543] = s[1] ? level0[1086] : level0[1087];
	assign level1[544] = s[1] ? level0[1088] : level0[1089];
	assign level1[545] = s[1] ? level0[1090] : level0[1091];
	assign level1[546] = s[1] ? level0[1092] : level0[1093];
	assign level1[547] = s[1] ? level0[1094] : level0[1095];
	assign level1[548] = s[1] ? level0[1096] : level0[1097];
	assign level1[549] = s[1] ? level0[1098] : level0[1099];
	assign level1[550] = s[1] ? level0[1100] : level0[1101];
	assign level1[551] = s[1] ? level0[1102] : level0[1103];
	assign level1[552] = s[1] ? level0[1104] : level0[1105];
	assign level1[553] = s[1] ? level0[1106] : level0[1107];
	assign level1[554] = s[1] ? level0[1108] : level0[1109];
	assign level1[555] = s[1] ? level0[1110] : level0[1111];
	assign level1[556] = s[1] ? level0[1112] : level0[1113];
	assign level1[557] = s[1] ? level0[1114] : level0[1115];
	assign level1[558] = s[1] ? level0[1116] : level0[1117];
	assign level1[559] = s[1] ? level0[1118] : level0[1119];
	assign level1[560] = s[1] ? level0[1120] : level0[1121];
	assign level1[561] = s[1] ? level0[1122] : level0[1123];
	assign level1[562] = s[1] ? level0[1124] : level0[1125];
	assign level1[563] = s[1] ? level0[1126] : level0[1127];
	assign level1[564] = s[1] ? level0[1128] : level0[1129];
	assign level1[565] = s[1] ? level0[1130] : level0[1131];
	assign level1[566] = s[1] ? level0[1132] : level0[1133];
	assign level1[567] = s[1] ? level0[1134] : level0[1135];
	assign level1[568] = s[1] ? level0[1136] : level0[1137];
	assign level1[569] = s[1] ? level0[1138] : level0[1139];
	assign level1[570] = s[1] ? level0[1140] : level0[1141];
	assign level1[571] = s[1] ? level0[1142] : level0[1143];
	assign level1[572] = s[1] ? level0[1144] : level0[1145];
	assign level1[573] = s[1] ? level0[1146] : level0[1147];
	assign level1[574] = s[1] ? level0[1148] : level0[1149];
	assign level1[575] = s[1] ? level0[1150] : level0[1151];
	assign level1[576] = s[1] ? level0[1152] : level0[1153];
	assign level1[577] = s[1] ? level0[1154] : level0[1155];
	assign level1[578] = s[1] ? level0[1156] : level0[1157];
	assign level1[579] = s[1] ? level0[1158] : level0[1159];
	assign level1[580] = s[1] ? level0[1160] : level0[1161];
	assign level1[581] = s[1] ? level0[1162] : level0[1163];
	assign level1[582] = s[1] ? level0[1164] : level0[1165];
	assign level1[583] = s[1] ? level0[1166] : level0[1167];
	assign level1[584] = s[1] ? level0[1168] : level0[1169];
	assign level1[585] = s[1] ? level0[1170] : level0[1171];
	assign level1[586] = s[1] ? level0[1172] : level0[1173];
	assign level1[587] = s[1] ? level0[1174] : level0[1175];
	assign level1[588] = s[1] ? level0[1176] : level0[1177];
	assign level1[589] = s[1] ? level0[1178] : level0[1179];
	assign level1[590] = s[1] ? level0[1180] : level0[1181];
	assign level1[591] = s[1] ? level0[1182] : level0[1183];
	assign level1[592] = s[1] ? level0[1184] : level0[1185];
	assign level1[593] = s[1] ? level0[1186] : level0[1187];
	assign level1[594] = s[1] ? level0[1188] : level0[1189];
	assign level1[595] = s[1] ? level0[1190] : level0[1191];
	assign level1[596] = s[1] ? level0[1192] : level0[1193];
	assign level1[597] = s[1] ? level0[1194] : level0[1195];
	assign level1[598] = s[1] ? level0[1196] : level0[1197];
	assign level1[599] = s[1] ? level0[1198] : level0[1199];
	assign level1[600] = s[1] ? level0[1200] : level0[1201];
	assign level1[601] = s[1] ? level0[1202] : level0[1203];
	assign level1[602] = s[1] ? level0[1204] : level0[1205];
	assign level1[603] = s[1] ? level0[1206] : level0[1207];
	assign level1[604] = s[1] ? level0[1208] : level0[1209];
	assign level1[605] = s[1] ? level0[1210] : level0[1211];
	assign level1[606] = s[1] ? level0[1212] : level0[1213];
	assign level1[607] = s[1] ? level0[1214] : level0[1215];
	assign level1[608] = s[1] ? level0[1216] : level0[1217];
	assign level1[609] = s[1] ? level0[1218] : level0[1219];
	assign level1[610] = s[1] ? level0[1220] : level0[1221];
	assign level1[611] = s[1] ? level0[1222] : level0[1223];
	assign level1[612] = s[1] ? level0[1224] : level0[1225];
	assign level1[613] = s[1] ? level0[1226] : level0[1227];
	assign level1[614] = s[1] ? level0[1228] : level0[1229];
	assign level1[615] = s[1] ? level0[1230] : level0[1231];
	assign level1[616] = s[1] ? level0[1232] : level0[1233];
	assign level1[617] = s[1] ? level0[1234] : level0[1235];
	assign level1[618] = s[1] ? level0[1236] : level0[1237];
	assign level1[619] = s[1] ? level0[1238] : level0[1239];
	assign level1[620] = s[1] ? level0[1240] : level0[1241];
	assign level1[621] = s[1] ? level0[1242] : level0[1243];
	assign level1[622] = s[1] ? level0[1244] : level0[1245];
	assign level1[623] = s[1] ? level0[1246] : level0[1247];
	assign level1[624] = s[1] ? level0[1248] : level0[1249];
	assign level1[625] = s[1] ? level0[1250] : level0[1251];
	assign level1[626] = s[1] ? level0[1252] : level0[1253];
	assign level1[627] = s[1] ? level0[1254] : level0[1255];
	assign level1[628] = s[1] ? level0[1256] : level0[1257];
	assign level1[629] = s[1] ? level0[1258] : level0[1259];
	assign level1[630] = s[1] ? level0[1260] : level0[1261];
	assign level1[631] = s[1] ? level0[1262] : level0[1263];
	assign level1[632] = s[1] ? level0[1264] : level0[1265];
	assign level1[633] = s[1] ? level0[1266] : level0[1267];
	assign level1[634] = s[1] ? level0[1268] : level0[1269];
	assign level1[635] = s[1] ? level0[1270] : level0[1271];
	assign level1[636] = s[1] ? level0[1272] : level0[1273];
	assign level1[637] = s[1] ? level0[1274] : level0[1275];
	assign level1[638] = s[1] ? level0[1276] : level0[1277];
	assign level1[639] = s[1] ? level0[1278] : level0[1279];
	assign level1[640] = s[1] ? level0[1280] : level0[1281];
	assign level1[641] = s[1] ? level0[1282] : level0[1283];
	assign level1[642] = s[1] ? level0[1284] : level0[1285];
	assign level1[643] = s[1] ? level0[1286] : level0[1287];
	assign level1[644] = s[1] ? level0[1288] : level0[1289];
	assign level1[645] = s[1] ? level0[1290] : level0[1291];
	assign level1[646] = s[1] ? level0[1292] : level0[1293];
	assign level1[647] = s[1] ? level0[1294] : level0[1295];
	assign level1[648] = s[1] ? level0[1296] : level0[1297];
	assign level1[649] = s[1] ? level0[1298] : level0[1299];
	assign level1[650] = s[1] ? level0[1300] : level0[1301];
	assign level1[651] = s[1] ? level0[1302] : level0[1303];
	assign level1[652] = s[1] ? level0[1304] : level0[1305];
	assign level1[653] = s[1] ? level0[1306] : level0[1307];
	assign level1[654] = s[1] ? level0[1308] : level0[1309];
	assign level1[655] = s[1] ? level0[1310] : level0[1311];
	assign level1[656] = s[1] ? level0[1312] : level0[1313];
	assign level1[657] = s[1] ? level0[1314] : level0[1315];
	assign level1[658] = s[1] ? level0[1316] : level0[1317];
	assign level1[659] = s[1] ? level0[1318] : level0[1319];
	assign level1[660] = s[1] ? level0[1320] : level0[1321];
	assign level1[661] = s[1] ? level0[1322] : level0[1323];
	assign level1[662] = s[1] ? level0[1324] : level0[1325];
	assign level1[663] = s[1] ? level0[1326] : level0[1327];
	assign level1[664] = s[1] ? level0[1328] : level0[1329];
	assign level1[665] = s[1] ? level0[1330] : level0[1331];
	assign level1[666] = s[1] ? level0[1332] : level0[1333];
	assign level1[667] = s[1] ? level0[1334] : level0[1335];
	assign level1[668] = s[1] ? level0[1336] : level0[1337];
	assign level1[669] = s[1] ? level0[1338] : level0[1339];
	assign level1[670] = s[1] ? level0[1340] : level0[1341];
	assign level1[671] = s[1] ? level0[1342] : level0[1343];
	assign level1[672] = s[1] ? level0[1344] : level0[1345];
	assign level1[673] = s[1] ? level0[1346] : level0[1347];
	assign level1[674] = s[1] ? level0[1348] : level0[1349];
	assign level1[675] = s[1] ? level0[1350] : level0[1351];
	assign level1[676] = s[1] ? level0[1352] : level0[1353];
	assign level1[677] = s[1] ? level0[1354] : level0[1355];
	assign level1[678] = s[1] ? level0[1356] : level0[1357];
	assign level1[679] = s[1] ? level0[1358] : level0[1359];
	assign level1[680] = s[1] ? level0[1360] : level0[1361];
	assign level1[681] = s[1] ? level0[1362] : level0[1363];
	assign level1[682] = s[1] ? level0[1364] : level0[1365];
	assign level1[683] = s[1] ? level0[1366] : level0[1367];
	assign level1[684] = s[1] ? level0[1368] : level0[1369];
	assign level1[685] = s[1] ? level0[1370] : level0[1371];
	assign level1[686] = s[1] ? level0[1372] : level0[1373];
	assign level1[687] = s[1] ? level0[1374] : level0[1375];
	assign level1[688] = s[1] ? level0[1376] : level0[1377];
	assign level1[689] = s[1] ? level0[1378] : level0[1379];
	assign level1[690] = s[1] ? level0[1380] : level0[1381];
	assign level1[691] = s[1] ? level0[1382] : level0[1383];
	assign level1[692] = s[1] ? level0[1384] : level0[1385];
	assign level1[693] = s[1] ? level0[1386] : level0[1387];
	assign level1[694] = s[1] ? level0[1388] : level0[1389];
	assign level1[695] = s[1] ? level0[1390] : level0[1391];
	assign level1[696] = s[1] ? level0[1392] : level0[1393];
	assign level1[697] = s[1] ? level0[1394] : level0[1395];
	assign level1[698] = s[1] ? level0[1396] : level0[1397];
	assign level1[699] = s[1] ? level0[1398] : level0[1399];
	assign level1[700] = s[1] ? level0[1400] : level0[1401];
	assign level1[701] = s[1] ? level0[1402] : level0[1403];
	assign level1[702] = s[1] ? level0[1404] : level0[1405];
	assign level1[703] = s[1] ? level0[1406] : level0[1407];
	assign level1[704] = s[1] ? level0[1408] : level0[1409];
	assign level1[705] = s[1] ? level0[1410] : level0[1411];
	assign level1[706] = s[1] ? level0[1412] : level0[1413];
	assign level1[707] = s[1] ? level0[1414] : level0[1415];
	assign level1[708] = s[1] ? level0[1416] : level0[1417];
	assign level1[709] = s[1] ? level0[1418] : level0[1419];
	assign level1[710] = s[1] ? level0[1420] : level0[1421];
	assign level1[711] = s[1] ? level0[1422] : level0[1423];
	assign level1[712] = s[1] ? level0[1424] : level0[1425];
	assign level1[713] = s[1] ? level0[1426] : level0[1427];
	assign level1[714] = s[1] ? level0[1428] : level0[1429];
	assign level1[715] = s[1] ? level0[1430] : level0[1431];
	assign level1[716] = s[1] ? level0[1432] : level0[1433];
	assign level1[717] = s[1] ? level0[1434] : level0[1435];
	assign level1[718] = s[1] ? level0[1436] : level0[1437];
	assign level1[719] = s[1] ? level0[1438] : level0[1439];
	assign level1[720] = s[1] ? level0[1440] : level0[1441];
	assign level1[721] = s[1] ? level0[1442] : level0[1443];
	assign level1[722] = s[1] ? level0[1444] : level0[1445];
	assign level1[723] = s[1] ? level0[1446] : level0[1447];
	assign level1[724] = s[1] ? level0[1448] : level0[1449];
	assign level1[725] = s[1] ? level0[1450] : level0[1451];
	assign level1[726] = s[1] ? level0[1452] : level0[1453];
	assign level1[727] = s[1] ? level0[1454] : level0[1455];
	assign level1[728] = s[1] ? level0[1456] : level0[1457];
	assign level1[729] = s[1] ? level0[1458] : level0[1459];
	assign level1[730] = s[1] ? level0[1460] : level0[1461];
	assign level1[731] = s[1] ? level0[1462] : level0[1463];
	assign level1[732] = s[1] ? level0[1464] : level0[1465];
	assign level1[733] = s[1] ? level0[1466] : level0[1467];
	assign level1[734] = s[1] ? level0[1468] : level0[1469];
	assign level1[735] = s[1] ? level0[1470] : level0[1471];
	assign level1[736] = s[1] ? level0[1472] : level0[1473];
	assign level1[737] = s[1] ? level0[1474] : level0[1475];
	assign level1[738] = s[1] ? level0[1476] : level0[1477];
	assign level1[739] = s[1] ? level0[1478] : level0[1479];
	assign level1[740] = s[1] ? level0[1480] : level0[1481];
	assign level1[741] = s[1] ? level0[1482] : level0[1483];
	assign level1[742] = s[1] ? level0[1484] : level0[1485];
	assign level1[743] = s[1] ? level0[1486] : level0[1487];
	assign level1[744] = s[1] ? level0[1488] : level0[1489];
	assign level1[745] = s[1] ? level0[1490] : level0[1491];
	assign level1[746] = s[1] ? level0[1492] : level0[1493];
	assign level1[747] = s[1] ? level0[1494] : level0[1495];
	assign level1[748] = s[1] ? level0[1496] : level0[1497];
	assign level1[749] = s[1] ? level0[1498] : level0[1499];
	assign level1[750] = s[1] ? level0[1500] : level0[1501];
	assign level1[751] = s[1] ? level0[1502] : level0[1503];
	assign level1[752] = s[1] ? level0[1504] : level0[1505];
	assign level1[753] = s[1] ? level0[1506] : level0[1507];
	assign level1[754] = s[1] ? level0[1508] : level0[1509];
	assign level1[755] = s[1] ? level0[1510] : level0[1511];
	assign level1[756] = s[1] ? level0[1512] : level0[1513];
	assign level1[757] = s[1] ? level0[1514] : level0[1515];
	assign level1[758] = s[1] ? level0[1516] : level0[1517];
	assign level1[759] = s[1] ? level0[1518] : level0[1519];
	assign level1[760] = s[1] ? level0[1520] : level0[1521];
	assign level1[761] = s[1] ? level0[1522] : level0[1523];
	assign level1[762] = s[1] ? level0[1524] : level0[1525];
	assign level1[763] = s[1] ? level0[1526] : level0[1527];
	assign level1[764] = s[1] ? level0[1528] : level0[1529];
	assign level1[765] = s[1] ? level0[1530] : level0[1531];
	assign level1[766] = s[1] ? level0[1532] : level0[1533];
	assign level1[767] = s[1] ? level0[1534] : level0[1535];
	assign level1[768] = s[1] ? level0[1536] : level0[1537];
	assign level1[769] = s[1] ? level0[1538] : level0[1539];
	assign level1[770] = s[1] ? level0[1540] : level0[1541];
	assign level1[771] = s[1] ? level0[1542] : level0[1543];
	assign level1[772] = s[1] ? level0[1544] : level0[1545];
	assign level1[773] = s[1] ? level0[1546] : level0[1547];
	assign level1[774] = s[1] ? level0[1548] : level0[1549];
	assign level1[775] = s[1] ? level0[1550] : level0[1551];
	assign level1[776] = s[1] ? level0[1552] : level0[1553];
	assign level1[777] = s[1] ? level0[1554] : level0[1555];
	assign level1[778] = s[1] ? level0[1556] : level0[1557];
	assign level1[779] = s[1] ? level0[1558] : level0[1559];
	assign level1[780] = s[1] ? level0[1560] : level0[1561];
	assign level1[781] = s[1] ? level0[1562] : level0[1563];
	assign level1[782] = s[1] ? level0[1564] : level0[1565];
	assign level1[783] = s[1] ? level0[1566] : level0[1567];
	assign level1[784] = s[1] ? level0[1568] : level0[1569];
	assign level1[785] = s[1] ? level0[1570] : level0[1571];
	assign level1[786] = s[1] ? level0[1572] : level0[1573];
	assign level1[787] = s[1] ? level0[1574] : level0[1575];
	assign level1[788] = s[1] ? level0[1576] : level0[1577];
	assign level1[789] = s[1] ? level0[1578] : level0[1579];
	assign level1[790] = s[1] ? level0[1580] : level0[1581];
	assign level1[791] = s[1] ? level0[1582] : level0[1583];
	assign level1[792] = s[1] ? level0[1584] : level0[1585];
	assign level1[793] = s[1] ? level0[1586] : level0[1587];
	assign level1[794] = s[1] ? level0[1588] : level0[1589];
	assign level1[795] = s[1] ? level0[1590] : level0[1591];
	assign level1[796] = s[1] ? level0[1592] : level0[1593];
	assign level1[797] = s[1] ? level0[1594] : level0[1595];
	assign level1[798] = s[1] ? level0[1596] : level0[1597];
	assign level1[799] = s[1] ? level0[1598] : level0[1599];
	assign level1[800] = s[1] ? level0[1600] : level0[1601];
	assign level1[801] = s[1] ? level0[1602] : level0[1603];
	assign level1[802] = s[1] ? level0[1604] : level0[1605];
	assign level1[803] = s[1] ? level0[1606] : level0[1607];
	assign level1[804] = s[1] ? level0[1608] : level0[1609];
	assign level1[805] = s[1] ? level0[1610] : level0[1611];
	assign level1[806] = s[1] ? level0[1612] : level0[1613];
	assign level1[807] = s[1] ? level0[1614] : level0[1615];
	assign level1[808] = s[1] ? level0[1616] : level0[1617];
	assign level1[809] = s[1] ? level0[1618] : level0[1619];
	assign level1[810] = s[1] ? level0[1620] : level0[1621];
	assign level1[811] = s[1] ? level0[1622] : level0[1623];
	assign level1[812] = s[1] ? level0[1624] : level0[1625];
	assign level1[813] = s[1] ? level0[1626] : level0[1627];
	assign level1[814] = s[1] ? level0[1628] : level0[1629];
	assign level1[815] = s[1] ? level0[1630] : level0[1631];
	assign level1[816] = s[1] ? level0[1632] : level0[1633];
	assign level1[817] = s[1] ? level0[1634] : level0[1635];
	assign level1[818] = s[1] ? level0[1636] : level0[1637];
	assign level1[819] = s[1] ? level0[1638] : level0[1639];
	assign level1[820] = s[1] ? level0[1640] : level0[1641];
	assign level1[821] = s[1] ? level0[1642] : level0[1643];
	assign level1[822] = s[1] ? level0[1644] : level0[1645];
	assign level1[823] = s[1] ? level0[1646] : level0[1647];
	assign level1[824] = s[1] ? level0[1648] : level0[1649];
	assign level1[825] = s[1] ? level0[1650] : level0[1651];
	assign level1[826] = s[1] ? level0[1652] : level0[1653];
	assign level1[827] = s[1] ? level0[1654] : level0[1655];
	assign level1[828] = s[1] ? level0[1656] : level0[1657];
	assign level1[829] = s[1] ? level0[1658] : level0[1659];
	assign level1[830] = s[1] ? level0[1660] : level0[1661];
	assign level1[831] = s[1] ? level0[1662] : level0[1663];
	assign level1[832] = s[1] ? level0[1664] : level0[1665];
	assign level1[833] = s[1] ? level0[1666] : level0[1667];
	assign level1[834] = s[1] ? level0[1668] : level0[1669];
	assign level1[835] = s[1] ? level0[1670] : level0[1671];
	assign level1[836] = s[1] ? level0[1672] : level0[1673];
	assign level1[837] = s[1] ? level0[1674] : level0[1675];
	assign level1[838] = s[1] ? level0[1676] : level0[1677];
	assign level1[839] = s[1] ? level0[1678] : level0[1679];
	assign level1[840] = s[1] ? level0[1680] : level0[1681];
	assign level1[841] = s[1] ? level0[1682] : level0[1683];
	assign level1[842] = s[1] ? level0[1684] : level0[1685];
	assign level1[843] = s[1] ? level0[1686] : level0[1687];
	assign level1[844] = s[1] ? level0[1688] : level0[1689];
	assign level1[845] = s[1] ? level0[1690] : level0[1691];
	assign level1[846] = s[1] ? level0[1692] : level0[1693];
	assign level1[847] = s[1] ? level0[1694] : level0[1695];
	assign level1[848] = s[1] ? level0[1696] : level0[1697];
	assign level1[849] = s[1] ? level0[1698] : level0[1699];
	assign level1[850] = s[1] ? level0[1700] : level0[1701];
	assign level1[851] = s[1] ? level0[1702] : level0[1703];
	assign level1[852] = s[1] ? level0[1704] : level0[1705];
	assign level1[853] = s[1] ? level0[1706] : level0[1707];
	assign level1[854] = s[1] ? level0[1708] : level0[1709];
	assign level1[855] = s[1] ? level0[1710] : level0[1711];
	assign level1[856] = s[1] ? level0[1712] : level0[1713];
	assign level1[857] = s[1] ? level0[1714] : level0[1715];
	assign level1[858] = s[1] ? level0[1716] : level0[1717];
	assign level1[859] = s[1] ? level0[1718] : level0[1719];
	assign level1[860] = s[1] ? level0[1720] : level0[1721];
	assign level1[861] = s[1] ? level0[1722] : level0[1723];
	assign level1[862] = s[1] ? level0[1724] : level0[1725];
	assign level1[863] = s[1] ? level0[1726] : level0[1727];
	assign level1[864] = s[1] ? level0[1728] : level0[1729];
	assign level1[865] = s[1] ? level0[1730] : level0[1731];
	assign level1[866] = s[1] ? level0[1732] : level0[1733];
	assign level1[867] = s[1] ? level0[1734] : level0[1735];
	assign level1[868] = s[1] ? level0[1736] : level0[1737];
	assign level1[869] = s[1] ? level0[1738] : level0[1739];
	assign level1[870] = s[1] ? level0[1740] : level0[1741];
	assign level1[871] = s[1] ? level0[1742] : level0[1743];
	assign level1[872] = s[1] ? level0[1744] : level0[1745];
	assign level1[873] = s[1] ? level0[1746] : level0[1747];
	assign level1[874] = s[1] ? level0[1748] : level0[1749];
	assign level1[875] = s[1] ? level0[1750] : level0[1751];
	assign level1[876] = s[1] ? level0[1752] : level0[1753];
	assign level1[877] = s[1] ? level0[1754] : level0[1755];
	assign level1[878] = s[1] ? level0[1756] : level0[1757];
	assign level1[879] = s[1] ? level0[1758] : level0[1759];
	assign level1[880] = s[1] ? level0[1760] : level0[1761];
	assign level1[881] = s[1] ? level0[1762] : level0[1763];
	assign level1[882] = s[1] ? level0[1764] : level0[1765];
	assign level1[883] = s[1] ? level0[1766] : level0[1767];
	assign level1[884] = s[1] ? level0[1768] : level0[1769];
	assign level1[885] = s[1] ? level0[1770] : level0[1771];
	assign level1[886] = s[1] ? level0[1772] : level0[1773];
	assign level1[887] = s[1] ? level0[1774] : level0[1775];
	assign level1[888] = s[1] ? level0[1776] : level0[1777];
	assign level1[889] = s[1] ? level0[1778] : level0[1779];
	assign level1[890] = s[1] ? level0[1780] : level0[1781];
	assign level1[891] = s[1] ? level0[1782] : level0[1783];
	assign level1[892] = s[1] ? level0[1784] : level0[1785];
	assign level1[893] = s[1] ? level0[1786] : level0[1787];
	assign level1[894] = s[1] ? level0[1788] : level0[1789];
	assign level1[895] = s[1] ? level0[1790] : level0[1791];
	assign level1[896] = s[1] ? level0[1792] : level0[1793];
	assign level1[897] = s[1] ? level0[1794] : level0[1795];
	assign level1[898] = s[1] ? level0[1796] : level0[1797];
	assign level1[899] = s[1] ? level0[1798] : level0[1799];
	assign level1[900] = s[1] ? level0[1800] : level0[1801];
	assign level1[901] = s[1] ? level0[1802] : level0[1803];
	assign level1[902] = s[1] ? level0[1804] : level0[1805];
	assign level1[903] = s[1] ? level0[1806] : level0[1807];
	assign level1[904] = s[1] ? level0[1808] : level0[1809];
	assign level1[905] = s[1] ? level0[1810] : level0[1811];
	assign level1[906] = s[1] ? level0[1812] : level0[1813];
	assign level1[907] = s[1] ? level0[1814] : level0[1815];
	assign level1[908] = s[1] ? level0[1816] : level0[1817];
	assign level1[909] = s[1] ? level0[1818] : level0[1819];
	assign level1[910] = s[1] ? level0[1820] : level0[1821];
	assign level1[911] = s[1] ? level0[1822] : level0[1823];
	assign level1[912] = s[1] ? level0[1824] : level0[1825];
	assign level1[913] = s[1] ? level0[1826] : level0[1827];
	assign level1[914] = s[1] ? level0[1828] : level0[1829];
	assign level1[915] = s[1] ? level0[1830] : level0[1831];
	assign level1[916] = s[1] ? level0[1832] : level0[1833];
	assign level1[917] = s[1] ? level0[1834] : level0[1835];
	assign level1[918] = s[1] ? level0[1836] : level0[1837];
	assign level1[919] = s[1] ? level0[1838] : level0[1839];
	assign level1[920] = s[1] ? level0[1840] : level0[1841];
	assign level1[921] = s[1] ? level0[1842] : level0[1843];
	assign level1[922] = s[1] ? level0[1844] : level0[1845];
	assign level1[923] = s[1] ? level0[1846] : level0[1847];
	assign level1[924] = s[1] ? level0[1848] : level0[1849];
	assign level1[925] = s[1] ? level0[1850] : level0[1851];
	assign level1[926] = s[1] ? level0[1852] : level0[1853];
	assign level1[927] = s[1] ? level0[1854] : level0[1855];
	assign level1[928] = s[1] ? level0[1856] : level0[1857];
	assign level1[929] = s[1] ? level0[1858] : level0[1859];
	assign level1[930] = s[1] ? level0[1860] : level0[1861];
	assign level1[931] = s[1] ? level0[1862] : level0[1863];
	assign level1[932] = s[1] ? level0[1864] : level0[1865];
	assign level1[933] = s[1] ? level0[1866] : level0[1867];
	assign level1[934] = s[1] ? level0[1868] : level0[1869];
	assign level1[935] = s[1] ? level0[1870] : level0[1871];
	assign level1[936] = s[1] ? level0[1872] : level0[1873];
	assign level1[937] = s[1] ? level0[1874] : level0[1875];
	assign level1[938] = s[1] ? level0[1876] : level0[1877];
	assign level1[939] = s[1] ? level0[1878] : level0[1879];
	assign level1[940] = s[1] ? level0[1880] : level0[1881];
	assign level1[941] = s[1] ? level0[1882] : level0[1883];
	assign level1[942] = s[1] ? level0[1884] : level0[1885];
	assign level1[943] = s[1] ? level0[1886] : level0[1887];
	assign level1[944] = s[1] ? level0[1888] : level0[1889];
	assign level1[945] = s[1] ? level0[1890] : level0[1891];
	assign level1[946] = s[1] ? level0[1892] : level0[1893];
	assign level1[947] = s[1] ? level0[1894] : level0[1895];
	assign level1[948] = s[1] ? level0[1896] : level0[1897];
	assign level1[949] = s[1] ? level0[1898] : level0[1899];
	assign level1[950] = s[1] ? level0[1900] : level0[1901];
	assign level1[951] = s[1] ? level0[1902] : level0[1903];
	assign level1[952] = s[1] ? level0[1904] : level0[1905];
	assign level1[953] = s[1] ? level0[1906] : level0[1907];
	assign level1[954] = s[1] ? level0[1908] : level0[1909];
	assign level1[955] = s[1] ? level0[1910] : level0[1911];
	assign level1[956] = s[1] ? level0[1912] : level0[1913];
	assign level1[957] = s[1] ? level0[1914] : level0[1915];
	assign level1[958] = s[1] ? level0[1916] : level0[1917];
	assign level1[959] = s[1] ? level0[1918] : level0[1919];
	assign level1[960] = s[1] ? level0[1920] : level0[1921];
	assign level1[961] = s[1] ? level0[1922] : level0[1923];
	assign level1[962] = s[1] ? level0[1924] : level0[1925];
	assign level1[963] = s[1] ? level0[1926] : level0[1927];
	assign level1[964] = s[1] ? level0[1928] : level0[1929];
	assign level1[965] = s[1] ? level0[1930] : level0[1931];
	assign level1[966] = s[1] ? level0[1932] : level0[1933];
	assign level1[967] = s[1] ? level0[1934] : level0[1935];
	assign level1[968] = s[1] ? level0[1936] : level0[1937];
	assign level1[969] = s[1] ? level0[1938] : level0[1939];
	assign level1[970] = s[1] ? level0[1940] : level0[1941];
	assign level1[971] = s[1] ? level0[1942] : level0[1943];
	assign level1[972] = s[1] ? level0[1944] : level0[1945];
	assign level1[973] = s[1] ? level0[1946] : level0[1947];
	assign level1[974] = s[1] ? level0[1948] : level0[1949];
	assign level1[975] = s[1] ? level0[1950] : level0[1951];
	assign level1[976] = s[1] ? level0[1952] : level0[1953];
	assign level1[977] = s[1] ? level0[1954] : level0[1955];
	assign level1[978] = s[1] ? level0[1956] : level0[1957];
	assign level1[979] = s[1] ? level0[1958] : level0[1959];
	assign level1[980] = s[1] ? level0[1960] : level0[1961];
	assign level1[981] = s[1] ? level0[1962] : level0[1963];
	assign level1[982] = s[1] ? level0[1964] : level0[1965];
	assign level1[983] = s[1] ? level0[1966] : level0[1967];
	assign level1[984] = s[1] ? level0[1968] : level0[1969];
	assign level1[985] = s[1] ? level0[1970] : level0[1971];
	assign level1[986] = s[1] ? level0[1972] : level0[1973];
	assign level1[987] = s[1] ? level0[1974] : level0[1975];
	assign level1[988] = s[1] ? level0[1976] : level0[1977];
	assign level1[989] = s[1] ? level0[1978] : level0[1979];
	assign level1[990] = s[1] ? level0[1980] : level0[1981];
	assign level1[991] = s[1] ? level0[1982] : level0[1983];
	assign level1[992] = s[1] ? level0[1984] : level0[1985];
	assign level1[993] = s[1] ? level0[1986] : level0[1987];
	assign level1[994] = s[1] ? level0[1988] : level0[1989];
	assign level1[995] = s[1] ? level0[1990] : level0[1991];
	assign level1[996] = s[1] ? level0[1992] : level0[1993];
	assign level1[997] = s[1] ? level0[1994] : level0[1995];
	assign level1[998] = s[1] ? level0[1996] : level0[1997];
	assign level1[999] = s[1] ? level0[1998] : level0[1999];
	assign level1[1000] = s[1] ? level0[2000] : level0[2001];
	assign level1[1001] = s[1] ? level0[2002] : level0[2003];
	assign level1[1002] = s[1] ? level0[2004] : level0[2005];
	assign level1[1003] = s[1] ? level0[2006] : level0[2007];
	assign level1[1004] = s[1] ? level0[2008] : level0[2009];
	assign level1[1005] = s[1] ? level0[2010] : level0[2011];
	assign level1[1006] = s[1] ? level0[2012] : level0[2013];
	assign level1[1007] = s[1] ? level0[2014] : level0[2015];
	assign level1[1008] = s[1] ? level0[2016] : level0[2017];
	assign level1[1009] = s[1] ? level0[2018] : level0[2019];
	assign level1[1010] = s[1] ? level0[2020] : level0[2021];
	assign level1[1011] = s[1] ? level0[2022] : level0[2023];
	assign level1[1012] = s[1] ? level0[2024] : level0[2025];
	assign level1[1013] = s[1] ? level0[2026] : level0[2027];
	assign level1[1014] = s[1] ? level0[2028] : level0[2029];
	assign level1[1015] = s[1] ? level0[2030] : level0[2031];
	assign level1[1016] = s[1] ? level0[2032] : level0[2033];
	assign level1[1017] = s[1] ? level0[2034] : level0[2035];
	assign level1[1018] = s[1] ? level0[2036] : level0[2037];
	assign level1[1019] = s[1] ? level0[2038] : level0[2039];
	assign level1[1020] = s[1] ? level0[2040] : level0[2041];
	assign level1[1021] = s[1] ? level0[2042] : level0[2043];
	assign level1[1022] = s[1] ? level0[2044] : level0[2045];
	assign level1[1023] = s[1] ? level0[2046] : level0[2047];

	assign level2[0] = s[2] ? level1[0] : level1[1];
	assign level2[1] = s[2] ? level1[2] : level1[3];
	assign level2[2] = s[2] ? level1[4] : level1[5];
	assign level2[3] = s[2] ? level1[6] : level1[7];
	assign level2[4] = s[2] ? level1[8] : level1[9];
	assign level2[5] = s[2] ? level1[10] : level1[11];
	assign level2[6] = s[2] ? level1[12] : level1[13];
	assign level2[7] = s[2] ? level1[14] : level1[15];
	assign level2[8] = s[2] ? level1[16] : level1[17];
	assign level2[9] = s[2] ? level1[18] : level1[19];
	assign level2[10] = s[2] ? level1[20] : level1[21];
	assign level2[11] = s[2] ? level1[22] : level1[23];
	assign level2[12] = s[2] ? level1[24] : level1[25];
	assign level2[13] = s[2] ? level1[26] : level1[27];
	assign level2[14] = s[2] ? level1[28] : level1[29];
	assign level2[15] = s[2] ? level1[30] : level1[31];
	assign level2[16] = s[2] ? level1[32] : level1[33];
	assign level2[17] = s[2] ? level1[34] : level1[35];
	assign level2[18] = s[2] ? level1[36] : level1[37];
	assign level2[19] = s[2] ? level1[38] : level1[39];
	assign level2[20] = s[2] ? level1[40] : level1[41];
	assign level2[21] = s[2] ? level1[42] : level1[43];
	assign level2[22] = s[2] ? level1[44] : level1[45];
	assign level2[23] = s[2] ? level1[46] : level1[47];
	assign level2[24] = s[2] ? level1[48] : level1[49];
	assign level2[25] = s[2] ? level1[50] : level1[51];
	assign level2[26] = s[2] ? level1[52] : level1[53];
	assign level2[27] = s[2] ? level1[54] : level1[55];
	assign level2[28] = s[2] ? level1[56] : level1[57];
	assign level2[29] = s[2] ? level1[58] : level1[59];
	assign level2[30] = s[2] ? level1[60] : level1[61];
	assign level2[31] = s[2] ? level1[62] : level1[63];
	assign level2[32] = s[2] ? level1[64] : level1[65];
	assign level2[33] = s[2] ? level1[66] : level1[67];
	assign level2[34] = s[2] ? level1[68] : level1[69];
	assign level2[35] = s[2] ? level1[70] : level1[71];
	assign level2[36] = s[2] ? level1[72] : level1[73];
	assign level2[37] = s[2] ? level1[74] : level1[75];
	assign level2[38] = s[2] ? level1[76] : level1[77];
	assign level2[39] = s[2] ? level1[78] : level1[79];
	assign level2[40] = s[2] ? level1[80] : level1[81];
	assign level2[41] = s[2] ? level1[82] : level1[83];
	assign level2[42] = s[2] ? level1[84] : level1[85];
	assign level2[43] = s[2] ? level1[86] : level1[87];
	assign level2[44] = s[2] ? level1[88] : level1[89];
	assign level2[45] = s[2] ? level1[90] : level1[91];
	assign level2[46] = s[2] ? level1[92] : level1[93];
	assign level2[47] = s[2] ? level1[94] : level1[95];
	assign level2[48] = s[2] ? level1[96] : level1[97];
	assign level2[49] = s[2] ? level1[98] : level1[99];
	assign level2[50] = s[2] ? level1[100] : level1[101];
	assign level2[51] = s[2] ? level1[102] : level1[103];
	assign level2[52] = s[2] ? level1[104] : level1[105];
	assign level2[53] = s[2] ? level1[106] : level1[107];
	assign level2[54] = s[2] ? level1[108] : level1[109];
	assign level2[55] = s[2] ? level1[110] : level1[111];
	assign level2[56] = s[2] ? level1[112] : level1[113];
	assign level2[57] = s[2] ? level1[114] : level1[115];
	assign level2[58] = s[2] ? level1[116] : level1[117];
	assign level2[59] = s[2] ? level1[118] : level1[119];
	assign level2[60] = s[2] ? level1[120] : level1[121];
	assign level2[61] = s[2] ? level1[122] : level1[123];
	assign level2[62] = s[2] ? level1[124] : level1[125];
	assign level2[63] = s[2] ? level1[126] : level1[127];
	assign level2[64] = s[2] ? level1[128] : level1[129];
	assign level2[65] = s[2] ? level1[130] : level1[131];
	assign level2[66] = s[2] ? level1[132] : level1[133];
	assign level2[67] = s[2] ? level1[134] : level1[135];
	assign level2[68] = s[2] ? level1[136] : level1[137];
	assign level2[69] = s[2] ? level1[138] : level1[139];
	assign level2[70] = s[2] ? level1[140] : level1[141];
	assign level2[71] = s[2] ? level1[142] : level1[143];
	assign level2[72] = s[2] ? level1[144] : level1[145];
	assign level2[73] = s[2] ? level1[146] : level1[147];
	assign level2[74] = s[2] ? level1[148] : level1[149];
	assign level2[75] = s[2] ? level1[150] : level1[151];
	assign level2[76] = s[2] ? level1[152] : level1[153];
	assign level2[77] = s[2] ? level1[154] : level1[155];
	assign level2[78] = s[2] ? level1[156] : level1[157];
	assign level2[79] = s[2] ? level1[158] : level1[159];
	assign level2[80] = s[2] ? level1[160] : level1[161];
	assign level2[81] = s[2] ? level1[162] : level1[163];
	assign level2[82] = s[2] ? level1[164] : level1[165];
	assign level2[83] = s[2] ? level1[166] : level1[167];
	assign level2[84] = s[2] ? level1[168] : level1[169];
	assign level2[85] = s[2] ? level1[170] : level1[171];
	assign level2[86] = s[2] ? level1[172] : level1[173];
	assign level2[87] = s[2] ? level1[174] : level1[175];
	assign level2[88] = s[2] ? level1[176] : level1[177];
	assign level2[89] = s[2] ? level1[178] : level1[179];
	assign level2[90] = s[2] ? level1[180] : level1[181];
	assign level2[91] = s[2] ? level1[182] : level1[183];
	assign level2[92] = s[2] ? level1[184] : level1[185];
	assign level2[93] = s[2] ? level1[186] : level1[187];
	assign level2[94] = s[2] ? level1[188] : level1[189];
	assign level2[95] = s[2] ? level1[190] : level1[191];
	assign level2[96] = s[2] ? level1[192] : level1[193];
	assign level2[97] = s[2] ? level1[194] : level1[195];
	assign level2[98] = s[2] ? level1[196] : level1[197];
	assign level2[99] = s[2] ? level1[198] : level1[199];
	assign level2[100] = s[2] ? level1[200] : level1[201];
	assign level2[101] = s[2] ? level1[202] : level1[203];
	assign level2[102] = s[2] ? level1[204] : level1[205];
	assign level2[103] = s[2] ? level1[206] : level1[207];
	assign level2[104] = s[2] ? level1[208] : level1[209];
	assign level2[105] = s[2] ? level1[210] : level1[211];
	assign level2[106] = s[2] ? level1[212] : level1[213];
	assign level2[107] = s[2] ? level1[214] : level1[215];
	assign level2[108] = s[2] ? level1[216] : level1[217];
	assign level2[109] = s[2] ? level1[218] : level1[219];
	assign level2[110] = s[2] ? level1[220] : level1[221];
	assign level2[111] = s[2] ? level1[222] : level1[223];
	assign level2[112] = s[2] ? level1[224] : level1[225];
	assign level2[113] = s[2] ? level1[226] : level1[227];
	assign level2[114] = s[2] ? level1[228] : level1[229];
	assign level2[115] = s[2] ? level1[230] : level1[231];
	assign level2[116] = s[2] ? level1[232] : level1[233];
	assign level2[117] = s[2] ? level1[234] : level1[235];
	assign level2[118] = s[2] ? level1[236] : level1[237];
	assign level2[119] = s[2] ? level1[238] : level1[239];
	assign level2[120] = s[2] ? level1[240] : level1[241];
	assign level2[121] = s[2] ? level1[242] : level1[243];
	assign level2[122] = s[2] ? level1[244] : level1[245];
	assign level2[123] = s[2] ? level1[246] : level1[247];
	assign level2[124] = s[2] ? level1[248] : level1[249];
	assign level2[125] = s[2] ? level1[250] : level1[251];
	assign level2[126] = s[2] ? level1[252] : level1[253];
	assign level2[127] = s[2] ? level1[254] : level1[255];
	assign level2[128] = s[2] ? level1[256] : level1[257];
	assign level2[129] = s[2] ? level1[258] : level1[259];
	assign level2[130] = s[2] ? level1[260] : level1[261];
	assign level2[131] = s[2] ? level1[262] : level1[263];
	assign level2[132] = s[2] ? level1[264] : level1[265];
	assign level2[133] = s[2] ? level1[266] : level1[267];
	assign level2[134] = s[2] ? level1[268] : level1[269];
	assign level2[135] = s[2] ? level1[270] : level1[271];
	assign level2[136] = s[2] ? level1[272] : level1[273];
	assign level2[137] = s[2] ? level1[274] : level1[275];
	assign level2[138] = s[2] ? level1[276] : level1[277];
	assign level2[139] = s[2] ? level1[278] : level1[279];
	assign level2[140] = s[2] ? level1[280] : level1[281];
	assign level2[141] = s[2] ? level1[282] : level1[283];
	assign level2[142] = s[2] ? level1[284] : level1[285];
	assign level2[143] = s[2] ? level1[286] : level1[287];
	assign level2[144] = s[2] ? level1[288] : level1[289];
	assign level2[145] = s[2] ? level1[290] : level1[291];
	assign level2[146] = s[2] ? level1[292] : level1[293];
	assign level2[147] = s[2] ? level1[294] : level1[295];
	assign level2[148] = s[2] ? level1[296] : level1[297];
	assign level2[149] = s[2] ? level1[298] : level1[299];
	assign level2[150] = s[2] ? level1[300] : level1[301];
	assign level2[151] = s[2] ? level1[302] : level1[303];
	assign level2[152] = s[2] ? level1[304] : level1[305];
	assign level2[153] = s[2] ? level1[306] : level1[307];
	assign level2[154] = s[2] ? level1[308] : level1[309];
	assign level2[155] = s[2] ? level1[310] : level1[311];
	assign level2[156] = s[2] ? level1[312] : level1[313];
	assign level2[157] = s[2] ? level1[314] : level1[315];
	assign level2[158] = s[2] ? level1[316] : level1[317];
	assign level2[159] = s[2] ? level1[318] : level1[319];
	assign level2[160] = s[2] ? level1[320] : level1[321];
	assign level2[161] = s[2] ? level1[322] : level1[323];
	assign level2[162] = s[2] ? level1[324] : level1[325];
	assign level2[163] = s[2] ? level1[326] : level1[327];
	assign level2[164] = s[2] ? level1[328] : level1[329];
	assign level2[165] = s[2] ? level1[330] : level1[331];
	assign level2[166] = s[2] ? level1[332] : level1[333];
	assign level2[167] = s[2] ? level1[334] : level1[335];
	assign level2[168] = s[2] ? level1[336] : level1[337];
	assign level2[169] = s[2] ? level1[338] : level1[339];
	assign level2[170] = s[2] ? level1[340] : level1[341];
	assign level2[171] = s[2] ? level1[342] : level1[343];
	assign level2[172] = s[2] ? level1[344] : level1[345];
	assign level2[173] = s[2] ? level1[346] : level1[347];
	assign level2[174] = s[2] ? level1[348] : level1[349];
	assign level2[175] = s[2] ? level1[350] : level1[351];
	assign level2[176] = s[2] ? level1[352] : level1[353];
	assign level2[177] = s[2] ? level1[354] : level1[355];
	assign level2[178] = s[2] ? level1[356] : level1[357];
	assign level2[179] = s[2] ? level1[358] : level1[359];
	assign level2[180] = s[2] ? level1[360] : level1[361];
	assign level2[181] = s[2] ? level1[362] : level1[363];
	assign level2[182] = s[2] ? level1[364] : level1[365];
	assign level2[183] = s[2] ? level1[366] : level1[367];
	assign level2[184] = s[2] ? level1[368] : level1[369];
	assign level2[185] = s[2] ? level1[370] : level1[371];
	assign level2[186] = s[2] ? level1[372] : level1[373];
	assign level2[187] = s[2] ? level1[374] : level1[375];
	assign level2[188] = s[2] ? level1[376] : level1[377];
	assign level2[189] = s[2] ? level1[378] : level1[379];
	assign level2[190] = s[2] ? level1[380] : level1[381];
	assign level2[191] = s[2] ? level1[382] : level1[383];
	assign level2[192] = s[2] ? level1[384] : level1[385];
	assign level2[193] = s[2] ? level1[386] : level1[387];
	assign level2[194] = s[2] ? level1[388] : level1[389];
	assign level2[195] = s[2] ? level1[390] : level1[391];
	assign level2[196] = s[2] ? level1[392] : level1[393];
	assign level2[197] = s[2] ? level1[394] : level1[395];
	assign level2[198] = s[2] ? level1[396] : level1[397];
	assign level2[199] = s[2] ? level1[398] : level1[399];
	assign level2[200] = s[2] ? level1[400] : level1[401];
	assign level2[201] = s[2] ? level1[402] : level1[403];
	assign level2[202] = s[2] ? level1[404] : level1[405];
	assign level2[203] = s[2] ? level1[406] : level1[407];
	assign level2[204] = s[2] ? level1[408] : level1[409];
	assign level2[205] = s[2] ? level1[410] : level1[411];
	assign level2[206] = s[2] ? level1[412] : level1[413];
	assign level2[207] = s[2] ? level1[414] : level1[415];
	assign level2[208] = s[2] ? level1[416] : level1[417];
	assign level2[209] = s[2] ? level1[418] : level1[419];
	assign level2[210] = s[2] ? level1[420] : level1[421];
	assign level2[211] = s[2] ? level1[422] : level1[423];
	assign level2[212] = s[2] ? level1[424] : level1[425];
	assign level2[213] = s[2] ? level1[426] : level1[427];
	assign level2[214] = s[2] ? level1[428] : level1[429];
	assign level2[215] = s[2] ? level1[430] : level1[431];
	assign level2[216] = s[2] ? level1[432] : level1[433];
	assign level2[217] = s[2] ? level1[434] : level1[435];
	assign level2[218] = s[2] ? level1[436] : level1[437];
	assign level2[219] = s[2] ? level1[438] : level1[439];
	assign level2[220] = s[2] ? level1[440] : level1[441];
	assign level2[221] = s[2] ? level1[442] : level1[443];
	assign level2[222] = s[2] ? level1[444] : level1[445];
	assign level2[223] = s[2] ? level1[446] : level1[447];
	assign level2[224] = s[2] ? level1[448] : level1[449];
	assign level2[225] = s[2] ? level1[450] : level1[451];
	assign level2[226] = s[2] ? level1[452] : level1[453];
	assign level2[227] = s[2] ? level1[454] : level1[455];
	assign level2[228] = s[2] ? level1[456] : level1[457];
	assign level2[229] = s[2] ? level1[458] : level1[459];
	assign level2[230] = s[2] ? level1[460] : level1[461];
	assign level2[231] = s[2] ? level1[462] : level1[463];
	assign level2[232] = s[2] ? level1[464] : level1[465];
	assign level2[233] = s[2] ? level1[466] : level1[467];
	assign level2[234] = s[2] ? level1[468] : level1[469];
	assign level2[235] = s[2] ? level1[470] : level1[471];
	assign level2[236] = s[2] ? level1[472] : level1[473];
	assign level2[237] = s[2] ? level1[474] : level1[475];
	assign level2[238] = s[2] ? level1[476] : level1[477];
	assign level2[239] = s[2] ? level1[478] : level1[479];
	assign level2[240] = s[2] ? level1[480] : level1[481];
	assign level2[241] = s[2] ? level1[482] : level1[483];
	assign level2[242] = s[2] ? level1[484] : level1[485];
	assign level2[243] = s[2] ? level1[486] : level1[487];
	assign level2[244] = s[2] ? level1[488] : level1[489];
	assign level2[245] = s[2] ? level1[490] : level1[491];
	assign level2[246] = s[2] ? level1[492] : level1[493];
	assign level2[247] = s[2] ? level1[494] : level1[495];
	assign level2[248] = s[2] ? level1[496] : level1[497];
	assign level2[249] = s[2] ? level1[498] : level1[499];
	assign level2[250] = s[2] ? level1[500] : level1[501];
	assign level2[251] = s[2] ? level1[502] : level1[503];
	assign level2[252] = s[2] ? level1[504] : level1[505];
	assign level2[253] = s[2] ? level1[506] : level1[507];
	assign level2[254] = s[2] ? level1[508] : level1[509];
	assign level2[255] = s[2] ? level1[510] : level1[511];
	assign level2[256] = s[2] ? level1[512] : level1[513];
	assign level2[257] = s[2] ? level1[514] : level1[515];
	assign level2[258] = s[2] ? level1[516] : level1[517];
	assign level2[259] = s[2] ? level1[518] : level1[519];
	assign level2[260] = s[2] ? level1[520] : level1[521];
	assign level2[261] = s[2] ? level1[522] : level1[523];
	assign level2[262] = s[2] ? level1[524] : level1[525];
	assign level2[263] = s[2] ? level1[526] : level1[527];
	assign level2[264] = s[2] ? level1[528] : level1[529];
	assign level2[265] = s[2] ? level1[530] : level1[531];
	assign level2[266] = s[2] ? level1[532] : level1[533];
	assign level2[267] = s[2] ? level1[534] : level1[535];
	assign level2[268] = s[2] ? level1[536] : level1[537];
	assign level2[269] = s[2] ? level1[538] : level1[539];
	assign level2[270] = s[2] ? level1[540] : level1[541];
	assign level2[271] = s[2] ? level1[542] : level1[543];
	assign level2[272] = s[2] ? level1[544] : level1[545];
	assign level2[273] = s[2] ? level1[546] : level1[547];
	assign level2[274] = s[2] ? level1[548] : level1[549];
	assign level2[275] = s[2] ? level1[550] : level1[551];
	assign level2[276] = s[2] ? level1[552] : level1[553];
	assign level2[277] = s[2] ? level1[554] : level1[555];
	assign level2[278] = s[2] ? level1[556] : level1[557];
	assign level2[279] = s[2] ? level1[558] : level1[559];
	assign level2[280] = s[2] ? level1[560] : level1[561];
	assign level2[281] = s[2] ? level1[562] : level1[563];
	assign level2[282] = s[2] ? level1[564] : level1[565];
	assign level2[283] = s[2] ? level1[566] : level1[567];
	assign level2[284] = s[2] ? level1[568] : level1[569];
	assign level2[285] = s[2] ? level1[570] : level1[571];
	assign level2[286] = s[2] ? level1[572] : level1[573];
	assign level2[287] = s[2] ? level1[574] : level1[575];
	assign level2[288] = s[2] ? level1[576] : level1[577];
	assign level2[289] = s[2] ? level1[578] : level1[579];
	assign level2[290] = s[2] ? level1[580] : level1[581];
	assign level2[291] = s[2] ? level1[582] : level1[583];
	assign level2[292] = s[2] ? level1[584] : level1[585];
	assign level2[293] = s[2] ? level1[586] : level1[587];
	assign level2[294] = s[2] ? level1[588] : level1[589];
	assign level2[295] = s[2] ? level1[590] : level1[591];
	assign level2[296] = s[2] ? level1[592] : level1[593];
	assign level2[297] = s[2] ? level1[594] : level1[595];
	assign level2[298] = s[2] ? level1[596] : level1[597];
	assign level2[299] = s[2] ? level1[598] : level1[599];
	assign level2[300] = s[2] ? level1[600] : level1[601];
	assign level2[301] = s[2] ? level1[602] : level1[603];
	assign level2[302] = s[2] ? level1[604] : level1[605];
	assign level2[303] = s[2] ? level1[606] : level1[607];
	assign level2[304] = s[2] ? level1[608] : level1[609];
	assign level2[305] = s[2] ? level1[610] : level1[611];
	assign level2[306] = s[2] ? level1[612] : level1[613];
	assign level2[307] = s[2] ? level1[614] : level1[615];
	assign level2[308] = s[2] ? level1[616] : level1[617];
	assign level2[309] = s[2] ? level1[618] : level1[619];
	assign level2[310] = s[2] ? level1[620] : level1[621];
	assign level2[311] = s[2] ? level1[622] : level1[623];
	assign level2[312] = s[2] ? level1[624] : level1[625];
	assign level2[313] = s[2] ? level1[626] : level1[627];
	assign level2[314] = s[2] ? level1[628] : level1[629];
	assign level2[315] = s[2] ? level1[630] : level1[631];
	assign level2[316] = s[2] ? level1[632] : level1[633];
	assign level2[317] = s[2] ? level1[634] : level1[635];
	assign level2[318] = s[2] ? level1[636] : level1[637];
	assign level2[319] = s[2] ? level1[638] : level1[639];
	assign level2[320] = s[2] ? level1[640] : level1[641];
	assign level2[321] = s[2] ? level1[642] : level1[643];
	assign level2[322] = s[2] ? level1[644] : level1[645];
	assign level2[323] = s[2] ? level1[646] : level1[647];
	assign level2[324] = s[2] ? level1[648] : level1[649];
	assign level2[325] = s[2] ? level1[650] : level1[651];
	assign level2[326] = s[2] ? level1[652] : level1[653];
	assign level2[327] = s[2] ? level1[654] : level1[655];
	assign level2[328] = s[2] ? level1[656] : level1[657];
	assign level2[329] = s[2] ? level1[658] : level1[659];
	assign level2[330] = s[2] ? level1[660] : level1[661];
	assign level2[331] = s[2] ? level1[662] : level1[663];
	assign level2[332] = s[2] ? level1[664] : level1[665];
	assign level2[333] = s[2] ? level1[666] : level1[667];
	assign level2[334] = s[2] ? level1[668] : level1[669];
	assign level2[335] = s[2] ? level1[670] : level1[671];
	assign level2[336] = s[2] ? level1[672] : level1[673];
	assign level2[337] = s[2] ? level1[674] : level1[675];
	assign level2[338] = s[2] ? level1[676] : level1[677];
	assign level2[339] = s[2] ? level1[678] : level1[679];
	assign level2[340] = s[2] ? level1[680] : level1[681];
	assign level2[341] = s[2] ? level1[682] : level1[683];
	assign level2[342] = s[2] ? level1[684] : level1[685];
	assign level2[343] = s[2] ? level1[686] : level1[687];
	assign level2[344] = s[2] ? level1[688] : level1[689];
	assign level2[345] = s[2] ? level1[690] : level1[691];
	assign level2[346] = s[2] ? level1[692] : level1[693];
	assign level2[347] = s[2] ? level1[694] : level1[695];
	assign level2[348] = s[2] ? level1[696] : level1[697];
	assign level2[349] = s[2] ? level1[698] : level1[699];
	assign level2[350] = s[2] ? level1[700] : level1[701];
	assign level2[351] = s[2] ? level1[702] : level1[703];
	assign level2[352] = s[2] ? level1[704] : level1[705];
	assign level2[353] = s[2] ? level1[706] : level1[707];
	assign level2[354] = s[2] ? level1[708] : level1[709];
	assign level2[355] = s[2] ? level1[710] : level1[711];
	assign level2[356] = s[2] ? level1[712] : level1[713];
	assign level2[357] = s[2] ? level1[714] : level1[715];
	assign level2[358] = s[2] ? level1[716] : level1[717];
	assign level2[359] = s[2] ? level1[718] : level1[719];
	assign level2[360] = s[2] ? level1[720] : level1[721];
	assign level2[361] = s[2] ? level1[722] : level1[723];
	assign level2[362] = s[2] ? level1[724] : level1[725];
	assign level2[363] = s[2] ? level1[726] : level1[727];
	assign level2[364] = s[2] ? level1[728] : level1[729];
	assign level2[365] = s[2] ? level1[730] : level1[731];
	assign level2[366] = s[2] ? level1[732] : level1[733];
	assign level2[367] = s[2] ? level1[734] : level1[735];
	assign level2[368] = s[2] ? level1[736] : level1[737];
	assign level2[369] = s[2] ? level1[738] : level1[739];
	assign level2[370] = s[2] ? level1[740] : level1[741];
	assign level2[371] = s[2] ? level1[742] : level1[743];
	assign level2[372] = s[2] ? level1[744] : level1[745];
	assign level2[373] = s[2] ? level1[746] : level1[747];
	assign level2[374] = s[2] ? level1[748] : level1[749];
	assign level2[375] = s[2] ? level1[750] : level1[751];
	assign level2[376] = s[2] ? level1[752] : level1[753];
	assign level2[377] = s[2] ? level1[754] : level1[755];
	assign level2[378] = s[2] ? level1[756] : level1[757];
	assign level2[379] = s[2] ? level1[758] : level1[759];
	assign level2[380] = s[2] ? level1[760] : level1[761];
	assign level2[381] = s[2] ? level1[762] : level1[763];
	assign level2[382] = s[2] ? level1[764] : level1[765];
	assign level2[383] = s[2] ? level1[766] : level1[767];
	assign level2[384] = s[2] ? level1[768] : level1[769];
	assign level2[385] = s[2] ? level1[770] : level1[771];
	assign level2[386] = s[2] ? level1[772] : level1[773];
	assign level2[387] = s[2] ? level1[774] : level1[775];
	assign level2[388] = s[2] ? level1[776] : level1[777];
	assign level2[389] = s[2] ? level1[778] : level1[779];
	assign level2[390] = s[2] ? level1[780] : level1[781];
	assign level2[391] = s[2] ? level1[782] : level1[783];
	assign level2[392] = s[2] ? level1[784] : level1[785];
	assign level2[393] = s[2] ? level1[786] : level1[787];
	assign level2[394] = s[2] ? level1[788] : level1[789];
	assign level2[395] = s[2] ? level1[790] : level1[791];
	assign level2[396] = s[2] ? level1[792] : level1[793];
	assign level2[397] = s[2] ? level1[794] : level1[795];
	assign level2[398] = s[2] ? level1[796] : level1[797];
	assign level2[399] = s[2] ? level1[798] : level1[799];
	assign level2[400] = s[2] ? level1[800] : level1[801];
	assign level2[401] = s[2] ? level1[802] : level1[803];
	assign level2[402] = s[2] ? level1[804] : level1[805];
	assign level2[403] = s[2] ? level1[806] : level1[807];
	assign level2[404] = s[2] ? level1[808] : level1[809];
	assign level2[405] = s[2] ? level1[810] : level1[811];
	assign level2[406] = s[2] ? level1[812] : level1[813];
	assign level2[407] = s[2] ? level1[814] : level1[815];
	assign level2[408] = s[2] ? level1[816] : level1[817];
	assign level2[409] = s[2] ? level1[818] : level1[819];
	assign level2[410] = s[2] ? level1[820] : level1[821];
	assign level2[411] = s[2] ? level1[822] : level1[823];
	assign level2[412] = s[2] ? level1[824] : level1[825];
	assign level2[413] = s[2] ? level1[826] : level1[827];
	assign level2[414] = s[2] ? level1[828] : level1[829];
	assign level2[415] = s[2] ? level1[830] : level1[831];
	assign level2[416] = s[2] ? level1[832] : level1[833];
	assign level2[417] = s[2] ? level1[834] : level1[835];
	assign level2[418] = s[2] ? level1[836] : level1[837];
	assign level2[419] = s[2] ? level1[838] : level1[839];
	assign level2[420] = s[2] ? level1[840] : level1[841];
	assign level2[421] = s[2] ? level1[842] : level1[843];
	assign level2[422] = s[2] ? level1[844] : level1[845];
	assign level2[423] = s[2] ? level1[846] : level1[847];
	assign level2[424] = s[2] ? level1[848] : level1[849];
	assign level2[425] = s[2] ? level1[850] : level1[851];
	assign level2[426] = s[2] ? level1[852] : level1[853];
	assign level2[427] = s[2] ? level1[854] : level1[855];
	assign level2[428] = s[2] ? level1[856] : level1[857];
	assign level2[429] = s[2] ? level1[858] : level1[859];
	assign level2[430] = s[2] ? level1[860] : level1[861];
	assign level2[431] = s[2] ? level1[862] : level1[863];
	assign level2[432] = s[2] ? level1[864] : level1[865];
	assign level2[433] = s[2] ? level1[866] : level1[867];
	assign level2[434] = s[2] ? level1[868] : level1[869];
	assign level2[435] = s[2] ? level1[870] : level1[871];
	assign level2[436] = s[2] ? level1[872] : level1[873];
	assign level2[437] = s[2] ? level1[874] : level1[875];
	assign level2[438] = s[2] ? level1[876] : level1[877];
	assign level2[439] = s[2] ? level1[878] : level1[879];
	assign level2[440] = s[2] ? level1[880] : level1[881];
	assign level2[441] = s[2] ? level1[882] : level1[883];
	assign level2[442] = s[2] ? level1[884] : level1[885];
	assign level2[443] = s[2] ? level1[886] : level1[887];
	assign level2[444] = s[2] ? level1[888] : level1[889];
	assign level2[445] = s[2] ? level1[890] : level1[891];
	assign level2[446] = s[2] ? level1[892] : level1[893];
	assign level2[447] = s[2] ? level1[894] : level1[895];
	assign level2[448] = s[2] ? level1[896] : level1[897];
	assign level2[449] = s[2] ? level1[898] : level1[899];
	assign level2[450] = s[2] ? level1[900] : level1[901];
	assign level2[451] = s[2] ? level1[902] : level1[903];
	assign level2[452] = s[2] ? level1[904] : level1[905];
	assign level2[453] = s[2] ? level1[906] : level1[907];
	assign level2[454] = s[2] ? level1[908] : level1[909];
	assign level2[455] = s[2] ? level1[910] : level1[911];
	assign level2[456] = s[2] ? level1[912] : level1[913];
	assign level2[457] = s[2] ? level1[914] : level1[915];
	assign level2[458] = s[2] ? level1[916] : level1[917];
	assign level2[459] = s[2] ? level1[918] : level1[919];
	assign level2[460] = s[2] ? level1[920] : level1[921];
	assign level2[461] = s[2] ? level1[922] : level1[923];
	assign level2[462] = s[2] ? level1[924] : level1[925];
	assign level2[463] = s[2] ? level1[926] : level1[927];
	assign level2[464] = s[2] ? level1[928] : level1[929];
	assign level2[465] = s[2] ? level1[930] : level1[931];
	assign level2[466] = s[2] ? level1[932] : level1[933];
	assign level2[467] = s[2] ? level1[934] : level1[935];
	assign level2[468] = s[2] ? level1[936] : level1[937];
	assign level2[469] = s[2] ? level1[938] : level1[939];
	assign level2[470] = s[2] ? level1[940] : level1[941];
	assign level2[471] = s[2] ? level1[942] : level1[943];
	assign level2[472] = s[2] ? level1[944] : level1[945];
	assign level2[473] = s[2] ? level1[946] : level1[947];
	assign level2[474] = s[2] ? level1[948] : level1[949];
	assign level2[475] = s[2] ? level1[950] : level1[951];
	assign level2[476] = s[2] ? level1[952] : level1[953];
	assign level2[477] = s[2] ? level1[954] : level1[955];
	assign level2[478] = s[2] ? level1[956] : level1[957];
	assign level2[479] = s[2] ? level1[958] : level1[959];
	assign level2[480] = s[2] ? level1[960] : level1[961];
	assign level2[481] = s[2] ? level1[962] : level1[963];
	assign level2[482] = s[2] ? level1[964] : level1[965];
	assign level2[483] = s[2] ? level1[966] : level1[967];
	assign level2[484] = s[2] ? level1[968] : level1[969];
	assign level2[485] = s[2] ? level1[970] : level1[971];
	assign level2[486] = s[2] ? level1[972] : level1[973];
	assign level2[487] = s[2] ? level1[974] : level1[975];
	assign level2[488] = s[2] ? level1[976] : level1[977];
	assign level2[489] = s[2] ? level1[978] : level1[979];
	assign level2[490] = s[2] ? level1[980] : level1[981];
	assign level2[491] = s[2] ? level1[982] : level1[983];
	assign level2[492] = s[2] ? level1[984] : level1[985];
	assign level2[493] = s[2] ? level1[986] : level1[987];
	assign level2[494] = s[2] ? level1[988] : level1[989];
	assign level2[495] = s[2] ? level1[990] : level1[991];
	assign level2[496] = s[2] ? level1[992] : level1[993];
	assign level2[497] = s[2] ? level1[994] : level1[995];
	assign level2[498] = s[2] ? level1[996] : level1[997];
	assign level2[499] = s[2] ? level1[998] : level1[999];
	assign level2[500] = s[2] ? level1[1000] : level1[1001];
	assign level2[501] = s[2] ? level1[1002] : level1[1003];
	assign level2[502] = s[2] ? level1[1004] : level1[1005];
	assign level2[503] = s[2] ? level1[1006] : level1[1007];
	assign level2[504] = s[2] ? level1[1008] : level1[1009];
	assign level2[505] = s[2] ? level1[1010] : level1[1011];
	assign level2[506] = s[2] ? level1[1012] : level1[1013];
	assign level2[507] = s[2] ? level1[1014] : level1[1015];
	assign level2[508] = s[2] ? level1[1016] : level1[1017];
	assign level2[509] = s[2] ? level1[1018] : level1[1019];
	assign level2[510] = s[2] ? level1[1020] : level1[1021];
	assign level2[511] = s[2] ? level1[1022] : level1[1023];

	assign level3[0] = s[3] ? level2[0] : level2[1];
	assign level3[1] = s[3] ? level2[2] : level2[3];
	assign level3[2] = s[3] ? level2[4] : level2[5];
	assign level3[3] = s[3] ? level2[6] : level2[7];
	assign level3[4] = s[3] ? level2[8] : level2[9];
	assign level3[5] = s[3] ? level2[10] : level2[11];
	assign level3[6] = s[3] ? level2[12] : level2[13];
	assign level3[7] = s[3] ? level2[14] : level2[15];
	assign level3[8] = s[3] ? level2[16] : level2[17];
	assign level3[9] = s[3] ? level2[18] : level2[19];
	assign level3[10] = s[3] ? level2[20] : level2[21];
	assign level3[11] = s[3] ? level2[22] : level2[23];
	assign level3[12] = s[3] ? level2[24] : level2[25];
	assign level3[13] = s[3] ? level2[26] : level2[27];
	assign level3[14] = s[3] ? level2[28] : level2[29];
	assign level3[15] = s[3] ? level2[30] : level2[31];
	assign level3[16] = s[3] ? level2[32] : level2[33];
	assign level3[17] = s[3] ? level2[34] : level2[35];
	assign level3[18] = s[3] ? level2[36] : level2[37];
	assign level3[19] = s[3] ? level2[38] : level2[39];
	assign level3[20] = s[3] ? level2[40] : level2[41];
	assign level3[21] = s[3] ? level2[42] : level2[43];
	assign level3[22] = s[3] ? level2[44] : level2[45];
	assign level3[23] = s[3] ? level2[46] : level2[47];
	assign level3[24] = s[3] ? level2[48] : level2[49];
	assign level3[25] = s[3] ? level2[50] : level2[51];
	assign level3[26] = s[3] ? level2[52] : level2[53];
	assign level3[27] = s[3] ? level2[54] : level2[55];
	assign level3[28] = s[3] ? level2[56] : level2[57];
	assign level3[29] = s[3] ? level2[58] : level2[59];
	assign level3[30] = s[3] ? level2[60] : level2[61];
	assign level3[31] = s[3] ? level2[62] : level2[63];
	assign level3[32] = s[3] ? level2[64] : level2[65];
	assign level3[33] = s[3] ? level2[66] : level2[67];
	assign level3[34] = s[3] ? level2[68] : level2[69];
	assign level3[35] = s[3] ? level2[70] : level2[71];
	assign level3[36] = s[3] ? level2[72] : level2[73];
	assign level3[37] = s[3] ? level2[74] : level2[75];
	assign level3[38] = s[3] ? level2[76] : level2[77];
	assign level3[39] = s[3] ? level2[78] : level2[79];
	assign level3[40] = s[3] ? level2[80] : level2[81];
	assign level3[41] = s[3] ? level2[82] : level2[83];
	assign level3[42] = s[3] ? level2[84] : level2[85];
	assign level3[43] = s[3] ? level2[86] : level2[87];
	assign level3[44] = s[3] ? level2[88] : level2[89];
	assign level3[45] = s[3] ? level2[90] : level2[91];
	assign level3[46] = s[3] ? level2[92] : level2[93];
	assign level3[47] = s[3] ? level2[94] : level2[95];
	assign level3[48] = s[3] ? level2[96] : level2[97];
	assign level3[49] = s[3] ? level2[98] : level2[99];
	assign level3[50] = s[3] ? level2[100] : level2[101];
	assign level3[51] = s[3] ? level2[102] : level2[103];
	assign level3[52] = s[3] ? level2[104] : level2[105];
	assign level3[53] = s[3] ? level2[106] : level2[107];
	assign level3[54] = s[3] ? level2[108] : level2[109];
	assign level3[55] = s[3] ? level2[110] : level2[111];
	assign level3[56] = s[3] ? level2[112] : level2[113];
	assign level3[57] = s[3] ? level2[114] : level2[115];
	assign level3[58] = s[3] ? level2[116] : level2[117];
	assign level3[59] = s[3] ? level2[118] : level2[119];
	assign level3[60] = s[3] ? level2[120] : level2[121];
	assign level3[61] = s[3] ? level2[122] : level2[123];
	assign level3[62] = s[3] ? level2[124] : level2[125];
	assign level3[63] = s[3] ? level2[126] : level2[127];
	assign level3[64] = s[3] ? level2[128] : level2[129];
	assign level3[65] = s[3] ? level2[130] : level2[131];
	assign level3[66] = s[3] ? level2[132] : level2[133];
	assign level3[67] = s[3] ? level2[134] : level2[135];
	assign level3[68] = s[3] ? level2[136] : level2[137];
	assign level3[69] = s[3] ? level2[138] : level2[139];
	assign level3[70] = s[3] ? level2[140] : level2[141];
	assign level3[71] = s[3] ? level2[142] : level2[143];
	assign level3[72] = s[3] ? level2[144] : level2[145];
	assign level3[73] = s[3] ? level2[146] : level2[147];
	assign level3[74] = s[3] ? level2[148] : level2[149];
	assign level3[75] = s[3] ? level2[150] : level2[151];
	assign level3[76] = s[3] ? level2[152] : level2[153];
	assign level3[77] = s[3] ? level2[154] : level2[155];
	assign level3[78] = s[3] ? level2[156] : level2[157];
	assign level3[79] = s[3] ? level2[158] : level2[159];
	assign level3[80] = s[3] ? level2[160] : level2[161];
	assign level3[81] = s[3] ? level2[162] : level2[163];
	assign level3[82] = s[3] ? level2[164] : level2[165];
	assign level3[83] = s[3] ? level2[166] : level2[167];
	assign level3[84] = s[3] ? level2[168] : level2[169];
	assign level3[85] = s[3] ? level2[170] : level2[171];
	assign level3[86] = s[3] ? level2[172] : level2[173];
	assign level3[87] = s[3] ? level2[174] : level2[175];
	assign level3[88] = s[3] ? level2[176] : level2[177];
	assign level3[89] = s[3] ? level2[178] : level2[179];
	assign level3[90] = s[3] ? level2[180] : level2[181];
	assign level3[91] = s[3] ? level2[182] : level2[183];
	assign level3[92] = s[3] ? level2[184] : level2[185];
	assign level3[93] = s[3] ? level2[186] : level2[187];
	assign level3[94] = s[3] ? level2[188] : level2[189];
	assign level3[95] = s[3] ? level2[190] : level2[191];
	assign level3[96] = s[3] ? level2[192] : level2[193];
	assign level3[97] = s[3] ? level2[194] : level2[195];
	assign level3[98] = s[3] ? level2[196] : level2[197];
	assign level3[99] = s[3] ? level2[198] : level2[199];
	assign level3[100] = s[3] ? level2[200] : level2[201];
	assign level3[101] = s[3] ? level2[202] : level2[203];
	assign level3[102] = s[3] ? level2[204] : level2[205];
	assign level3[103] = s[3] ? level2[206] : level2[207];
	assign level3[104] = s[3] ? level2[208] : level2[209];
	assign level3[105] = s[3] ? level2[210] : level2[211];
	assign level3[106] = s[3] ? level2[212] : level2[213];
	assign level3[107] = s[3] ? level2[214] : level2[215];
	assign level3[108] = s[3] ? level2[216] : level2[217];
	assign level3[109] = s[3] ? level2[218] : level2[219];
	assign level3[110] = s[3] ? level2[220] : level2[221];
	assign level3[111] = s[3] ? level2[222] : level2[223];
	assign level3[112] = s[3] ? level2[224] : level2[225];
	assign level3[113] = s[3] ? level2[226] : level2[227];
	assign level3[114] = s[3] ? level2[228] : level2[229];
	assign level3[115] = s[3] ? level2[230] : level2[231];
	assign level3[116] = s[3] ? level2[232] : level2[233];
	assign level3[117] = s[3] ? level2[234] : level2[235];
	assign level3[118] = s[3] ? level2[236] : level2[237];
	assign level3[119] = s[3] ? level2[238] : level2[239];
	assign level3[120] = s[3] ? level2[240] : level2[241];
	assign level3[121] = s[3] ? level2[242] : level2[243];
	assign level3[122] = s[3] ? level2[244] : level2[245];
	assign level3[123] = s[3] ? level2[246] : level2[247];
	assign level3[124] = s[3] ? level2[248] : level2[249];
	assign level3[125] = s[3] ? level2[250] : level2[251];
	assign level3[126] = s[3] ? level2[252] : level2[253];
	assign level3[127] = s[3] ? level2[254] : level2[255];
	assign level3[128] = s[3] ? level2[256] : level2[257];
	assign level3[129] = s[3] ? level2[258] : level2[259];
	assign level3[130] = s[3] ? level2[260] : level2[261];
	assign level3[131] = s[3] ? level2[262] : level2[263];
	assign level3[132] = s[3] ? level2[264] : level2[265];
	assign level3[133] = s[3] ? level2[266] : level2[267];
	assign level3[134] = s[3] ? level2[268] : level2[269];
	assign level3[135] = s[3] ? level2[270] : level2[271];
	assign level3[136] = s[3] ? level2[272] : level2[273];
	assign level3[137] = s[3] ? level2[274] : level2[275];
	assign level3[138] = s[3] ? level2[276] : level2[277];
	assign level3[139] = s[3] ? level2[278] : level2[279];
	assign level3[140] = s[3] ? level2[280] : level2[281];
	assign level3[141] = s[3] ? level2[282] : level2[283];
	assign level3[142] = s[3] ? level2[284] : level2[285];
	assign level3[143] = s[3] ? level2[286] : level2[287];
	assign level3[144] = s[3] ? level2[288] : level2[289];
	assign level3[145] = s[3] ? level2[290] : level2[291];
	assign level3[146] = s[3] ? level2[292] : level2[293];
	assign level3[147] = s[3] ? level2[294] : level2[295];
	assign level3[148] = s[3] ? level2[296] : level2[297];
	assign level3[149] = s[3] ? level2[298] : level2[299];
	assign level3[150] = s[3] ? level2[300] : level2[301];
	assign level3[151] = s[3] ? level2[302] : level2[303];
	assign level3[152] = s[3] ? level2[304] : level2[305];
	assign level3[153] = s[3] ? level2[306] : level2[307];
	assign level3[154] = s[3] ? level2[308] : level2[309];
	assign level3[155] = s[3] ? level2[310] : level2[311];
	assign level3[156] = s[3] ? level2[312] : level2[313];
	assign level3[157] = s[3] ? level2[314] : level2[315];
	assign level3[158] = s[3] ? level2[316] : level2[317];
	assign level3[159] = s[3] ? level2[318] : level2[319];
	assign level3[160] = s[3] ? level2[320] : level2[321];
	assign level3[161] = s[3] ? level2[322] : level2[323];
	assign level3[162] = s[3] ? level2[324] : level2[325];
	assign level3[163] = s[3] ? level2[326] : level2[327];
	assign level3[164] = s[3] ? level2[328] : level2[329];
	assign level3[165] = s[3] ? level2[330] : level2[331];
	assign level3[166] = s[3] ? level2[332] : level2[333];
	assign level3[167] = s[3] ? level2[334] : level2[335];
	assign level3[168] = s[3] ? level2[336] : level2[337];
	assign level3[169] = s[3] ? level2[338] : level2[339];
	assign level3[170] = s[3] ? level2[340] : level2[341];
	assign level3[171] = s[3] ? level2[342] : level2[343];
	assign level3[172] = s[3] ? level2[344] : level2[345];
	assign level3[173] = s[3] ? level2[346] : level2[347];
	assign level3[174] = s[3] ? level2[348] : level2[349];
	assign level3[175] = s[3] ? level2[350] : level2[351];
	assign level3[176] = s[3] ? level2[352] : level2[353];
	assign level3[177] = s[3] ? level2[354] : level2[355];
	assign level3[178] = s[3] ? level2[356] : level2[357];
	assign level3[179] = s[3] ? level2[358] : level2[359];
	assign level3[180] = s[3] ? level2[360] : level2[361];
	assign level3[181] = s[3] ? level2[362] : level2[363];
	assign level3[182] = s[3] ? level2[364] : level2[365];
	assign level3[183] = s[3] ? level2[366] : level2[367];
	assign level3[184] = s[3] ? level2[368] : level2[369];
	assign level3[185] = s[3] ? level2[370] : level2[371];
	assign level3[186] = s[3] ? level2[372] : level2[373];
	assign level3[187] = s[3] ? level2[374] : level2[375];
	assign level3[188] = s[3] ? level2[376] : level2[377];
	assign level3[189] = s[3] ? level2[378] : level2[379];
	assign level3[190] = s[3] ? level2[380] : level2[381];
	assign level3[191] = s[3] ? level2[382] : level2[383];
	assign level3[192] = s[3] ? level2[384] : level2[385];
	assign level3[193] = s[3] ? level2[386] : level2[387];
	assign level3[194] = s[3] ? level2[388] : level2[389];
	assign level3[195] = s[3] ? level2[390] : level2[391];
	assign level3[196] = s[3] ? level2[392] : level2[393];
	assign level3[197] = s[3] ? level2[394] : level2[395];
	assign level3[198] = s[3] ? level2[396] : level2[397];
	assign level3[199] = s[3] ? level2[398] : level2[399];
	assign level3[200] = s[3] ? level2[400] : level2[401];
	assign level3[201] = s[3] ? level2[402] : level2[403];
	assign level3[202] = s[3] ? level2[404] : level2[405];
	assign level3[203] = s[3] ? level2[406] : level2[407];
	assign level3[204] = s[3] ? level2[408] : level2[409];
	assign level3[205] = s[3] ? level2[410] : level2[411];
	assign level3[206] = s[3] ? level2[412] : level2[413];
	assign level3[207] = s[3] ? level2[414] : level2[415];
	assign level3[208] = s[3] ? level2[416] : level2[417];
	assign level3[209] = s[3] ? level2[418] : level2[419];
	assign level3[210] = s[3] ? level2[420] : level2[421];
	assign level3[211] = s[3] ? level2[422] : level2[423];
	assign level3[212] = s[3] ? level2[424] : level2[425];
	assign level3[213] = s[3] ? level2[426] : level2[427];
	assign level3[214] = s[3] ? level2[428] : level2[429];
	assign level3[215] = s[3] ? level2[430] : level2[431];
	assign level3[216] = s[3] ? level2[432] : level2[433];
	assign level3[217] = s[3] ? level2[434] : level2[435];
	assign level3[218] = s[3] ? level2[436] : level2[437];
	assign level3[219] = s[3] ? level2[438] : level2[439];
	assign level3[220] = s[3] ? level2[440] : level2[441];
	assign level3[221] = s[3] ? level2[442] : level2[443];
	assign level3[222] = s[3] ? level2[444] : level2[445];
	assign level3[223] = s[3] ? level2[446] : level2[447];
	assign level3[224] = s[3] ? level2[448] : level2[449];
	assign level3[225] = s[3] ? level2[450] : level2[451];
	assign level3[226] = s[3] ? level2[452] : level2[453];
	assign level3[227] = s[3] ? level2[454] : level2[455];
	assign level3[228] = s[3] ? level2[456] : level2[457];
	assign level3[229] = s[3] ? level2[458] : level2[459];
	assign level3[230] = s[3] ? level2[460] : level2[461];
	assign level3[231] = s[3] ? level2[462] : level2[463];
	assign level3[232] = s[3] ? level2[464] : level2[465];
	assign level3[233] = s[3] ? level2[466] : level2[467];
	assign level3[234] = s[3] ? level2[468] : level2[469];
	assign level3[235] = s[3] ? level2[470] : level2[471];
	assign level3[236] = s[3] ? level2[472] : level2[473];
	assign level3[237] = s[3] ? level2[474] : level2[475];
	assign level3[238] = s[3] ? level2[476] : level2[477];
	assign level3[239] = s[3] ? level2[478] : level2[479];
	assign level3[240] = s[3] ? level2[480] : level2[481];
	assign level3[241] = s[3] ? level2[482] : level2[483];
	assign level3[242] = s[3] ? level2[484] : level2[485];
	assign level3[243] = s[3] ? level2[486] : level2[487];
	assign level3[244] = s[3] ? level2[488] : level2[489];
	assign level3[245] = s[3] ? level2[490] : level2[491];
	assign level3[246] = s[3] ? level2[492] : level2[493];
	assign level3[247] = s[3] ? level2[494] : level2[495];
	assign level3[248] = s[3] ? level2[496] : level2[497];
	assign level3[249] = s[3] ? level2[498] : level2[499];
	assign level3[250] = s[3] ? level2[500] : level2[501];
	assign level3[251] = s[3] ? level2[502] : level2[503];
	assign level3[252] = s[3] ? level2[504] : level2[505];
	assign level3[253] = s[3] ? level2[506] : level2[507];
	assign level3[254] = s[3] ? level2[508] : level2[509];
	assign level3[255] = s[3] ? level2[510] : level2[511];

	assign level4[0] = s[4] ? level3[0] : level3[1];
	assign level4[1] = s[4] ? level3[2] : level3[3];
	assign level4[2] = s[4] ? level3[4] : level3[5];
	assign level4[3] = s[4] ? level3[6] : level3[7];
	assign level4[4] = s[4] ? level3[8] : level3[9];
	assign level4[5] = s[4] ? level3[10] : level3[11];
	assign level4[6] = s[4] ? level3[12] : level3[13];
	assign level4[7] = s[4] ? level3[14] : level3[15];
	assign level4[8] = s[4] ? level3[16] : level3[17];
	assign level4[9] = s[4] ? level3[18] : level3[19];
	assign level4[10] = s[4] ? level3[20] : level3[21];
	assign level4[11] = s[4] ? level3[22] : level3[23];
	assign level4[12] = s[4] ? level3[24] : level3[25];
	assign level4[13] = s[4] ? level3[26] : level3[27];
	assign level4[14] = s[4] ? level3[28] : level3[29];
	assign level4[15] = s[4] ? level3[30] : level3[31];
	assign level4[16] = s[4] ? level3[32] : level3[33];
	assign level4[17] = s[4] ? level3[34] : level3[35];
	assign level4[18] = s[4] ? level3[36] : level3[37];
	assign level4[19] = s[4] ? level3[38] : level3[39];
	assign level4[20] = s[4] ? level3[40] : level3[41];
	assign level4[21] = s[4] ? level3[42] : level3[43];
	assign level4[22] = s[4] ? level3[44] : level3[45];
	assign level4[23] = s[4] ? level3[46] : level3[47];
	assign level4[24] = s[4] ? level3[48] : level3[49];
	assign level4[25] = s[4] ? level3[50] : level3[51];
	assign level4[26] = s[4] ? level3[52] : level3[53];
	assign level4[27] = s[4] ? level3[54] : level3[55];
	assign level4[28] = s[4] ? level3[56] : level3[57];
	assign level4[29] = s[4] ? level3[58] : level3[59];
	assign level4[30] = s[4] ? level3[60] : level3[61];
	assign level4[31] = s[4] ? level3[62] : level3[63];
	assign level4[32] = s[4] ? level3[64] : level3[65];
	assign level4[33] = s[4] ? level3[66] : level3[67];
	assign level4[34] = s[4] ? level3[68] : level3[69];
	assign level4[35] = s[4] ? level3[70] : level3[71];
	assign level4[36] = s[4] ? level3[72] : level3[73];
	assign level4[37] = s[4] ? level3[74] : level3[75];
	assign level4[38] = s[4] ? level3[76] : level3[77];
	assign level4[39] = s[4] ? level3[78] : level3[79];
	assign level4[40] = s[4] ? level3[80] : level3[81];
	assign level4[41] = s[4] ? level3[82] : level3[83];
	assign level4[42] = s[4] ? level3[84] : level3[85];
	assign level4[43] = s[4] ? level3[86] : level3[87];
	assign level4[44] = s[4] ? level3[88] : level3[89];
	assign level4[45] = s[4] ? level3[90] : level3[91];
	assign level4[46] = s[4] ? level3[92] : level3[93];
	assign level4[47] = s[4] ? level3[94] : level3[95];
	assign level4[48] = s[4] ? level3[96] : level3[97];
	assign level4[49] = s[4] ? level3[98] : level3[99];
	assign level4[50] = s[4] ? level3[100] : level3[101];
	assign level4[51] = s[4] ? level3[102] : level3[103];
	assign level4[52] = s[4] ? level3[104] : level3[105];
	assign level4[53] = s[4] ? level3[106] : level3[107];
	assign level4[54] = s[4] ? level3[108] : level3[109];
	assign level4[55] = s[4] ? level3[110] : level3[111];
	assign level4[56] = s[4] ? level3[112] : level3[113];
	assign level4[57] = s[4] ? level3[114] : level3[115];
	assign level4[58] = s[4] ? level3[116] : level3[117];
	assign level4[59] = s[4] ? level3[118] : level3[119];
	assign level4[60] = s[4] ? level3[120] : level3[121];
	assign level4[61] = s[4] ? level3[122] : level3[123];
	assign level4[62] = s[4] ? level3[124] : level3[125];
	assign level4[63] = s[4] ? level3[126] : level3[127];
	assign level4[64] = s[4] ? level3[128] : level3[129];
	assign level4[65] = s[4] ? level3[130] : level3[131];
	assign level4[66] = s[4] ? level3[132] : level3[133];
	assign level4[67] = s[4] ? level3[134] : level3[135];
	assign level4[68] = s[4] ? level3[136] : level3[137];
	assign level4[69] = s[4] ? level3[138] : level3[139];
	assign level4[70] = s[4] ? level3[140] : level3[141];
	assign level4[71] = s[4] ? level3[142] : level3[143];
	assign level4[72] = s[4] ? level3[144] : level3[145];
	assign level4[73] = s[4] ? level3[146] : level3[147];
	assign level4[74] = s[4] ? level3[148] : level3[149];
	assign level4[75] = s[4] ? level3[150] : level3[151];
	assign level4[76] = s[4] ? level3[152] : level3[153];
	assign level4[77] = s[4] ? level3[154] : level3[155];
	assign level4[78] = s[4] ? level3[156] : level3[157];
	assign level4[79] = s[4] ? level3[158] : level3[159];
	assign level4[80] = s[4] ? level3[160] : level3[161];
	assign level4[81] = s[4] ? level3[162] : level3[163];
	assign level4[82] = s[4] ? level3[164] : level3[165];
	assign level4[83] = s[4] ? level3[166] : level3[167];
	assign level4[84] = s[4] ? level3[168] : level3[169];
	assign level4[85] = s[4] ? level3[170] : level3[171];
	assign level4[86] = s[4] ? level3[172] : level3[173];
	assign level4[87] = s[4] ? level3[174] : level3[175];
	assign level4[88] = s[4] ? level3[176] : level3[177];
	assign level4[89] = s[4] ? level3[178] : level3[179];
	assign level4[90] = s[4] ? level3[180] : level3[181];
	assign level4[91] = s[4] ? level3[182] : level3[183];
	assign level4[92] = s[4] ? level3[184] : level3[185];
	assign level4[93] = s[4] ? level3[186] : level3[187];
	assign level4[94] = s[4] ? level3[188] : level3[189];
	assign level4[95] = s[4] ? level3[190] : level3[191];
	assign level4[96] = s[4] ? level3[192] : level3[193];
	assign level4[97] = s[4] ? level3[194] : level3[195];
	assign level4[98] = s[4] ? level3[196] : level3[197];
	assign level4[99] = s[4] ? level3[198] : level3[199];
	assign level4[100] = s[4] ? level3[200] : level3[201];
	assign level4[101] = s[4] ? level3[202] : level3[203];
	assign level4[102] = s[4] ? level3[204] : level3[205];
	assign level4[103] = s[4] ? level3[206] : level3[207];
	assign level4[104] = s[4] ? level3[208] : level3[209];
	assign level4[105] = s[4] ? level3[210] : level3[211];
	assign level4[106] = s[4] ? level3[212] : level3[213];
	assign level4[107] = s[4] ? level3[214] : level3[215];
	assign level4[108] = s[4] ? level3[216] : level3[217];
	assign level4[109] = s[4] ? level3[218] : level3[219];
	assign level4[110] = s[4] ? level3[220] : level3[221];
	assign level4[111] = s[4] ? level3[222] : level3[223];
	assign level4[112] = s[4] ? level3[224] : level3[225];
	assign level4[113] = s[4] ? level3[226] : level3[227];
	assign level4[114] = s[4] ? level3[228] : level3[229];
	assign level4[115] = s[4] ? level3[230] : level3[231];
	assign level4[116] = s[4] ? level3[232] : level3[233];
	assign level4[117] = s[4] ? level3[234] : level3[235];
	assign level4[118] = s[4] ? level3[236] : level3[237];
	assign level4[119] = s[4] ? level3[238] : level3[239];
	assign level4[120] = s[4] ? level3[240] : level3[241];
	assign level4[121] = s[4] ? level3[242] : level3[243];
	assign level4[122] = s[4] ? level3[244] : level3[245];
	assign level4[123] = s[4] ? level3[246] : level3[247];
	assign level4[124] = s[4] ? level3[248] : level3[249];
	assign level4[125] = s[4] ? level3[250] : level3[251];
	assign level4[126] = s[4] ? level3[252] : level3[253];
	assign level4[127] = s[4] ? level3[254] : level3[255];

	assign level5[0] = s[5] ? level4[0] : level4[1];
	assign level5[1] = s[5] ? level4[2] : level4[3];
	assign level5[2] = s[5] ? level4[4] : level4[5];
	assign level5[3] = s[5] ? level4[6] : level4[7];
	assign level5[4] = s[5] ? level4[8] : level4[9];
	assign level5[5] = s[5] ? level4[10] : level4[11];
	assign level5[6] = s[5] ? level4[12] : level4[13];
	assign level5[7] = s[5] ? level4[14] : level4[15];
	assign level5[8] = s[5] ? level4[16] : level4[17];
	assign level5[9] = s[5] ? level4[18] : level4[19];
	assign level5[10] = s[5] ? level4[20] : level4[21];
	assign level5[11] = s[5] ? level4[22] : level4[23];
	assign level5[12] = s[5] ? level4[24] : level4[25];
	assign level5[13] = s[5] ? level4[26] : level4[27];
	assign level5[14] = s[5] ? level4[28] : level4[29];
	assign level5[15] = s[5] ? level4[30] : level4[31];
	assign level5[16] = s[5] ? level4[32] : level4[33];
	assign level5[17] = s[5] ? level4[34] : level4[35];
	assign level5[18] = s[5] ? level4[36] : level4[37];
	assign level5[19] = s[5] ? level4[38] : level4[39];
	assign level5[20] = s[5] ? level4[40] : level4[41];
	assign level5[21] = s[5] ? level4[42] : level4[43];
	assign level5[22] = s[5] ? level4[44] : level4[45];
	assign level5[23] = s[5] ? level4[46] : level4[47];
	assign level5[24] = s[5] ? level4[48] : level4[49];
	assign level5[25] = s[5] ? level4[50] : level4[51];
	assign level5[26] = s[5] ? level4[52] : level4[53];
	assign level5[27] = s[5] ? level4[54] : level4[55];
	assign level5[28] = s[5] ? level4[56] : level4[57];
	assign level5[29] = s[5] ? level4[58] : level4[59];
	assign level5[30] = s[5] ? level4[60] : level4[61];
	assign level5[31] = s[5] ? level4[62] : level4[63];
	assign level5[32] = s[5] ? level4[64] : level4[65];
	assign level5[33] = s[5] ? level4[66] : level4[67];
	assign level5[34] = s[5] ? level4[68] : level4[69];
	assign level5[35] = s[5] ? level4[70] : level4[71];
	assign level5[36] = s[5] ? level4[72] : level4[73];
	assign level5[37] = s[5] ? level4[74] : level4[75];
	assign level5[38] = s[5] ? level4[76] : level4[77];
	assign level5[39] = s[5] ? level4[78] : level4[79];
	assign level5[40] = s[5] ? level4[80] : level4[81];
	assign level5[41] = s[5] ? level4[82] : level4[83];
	assign level5[42] = s[5] ? level4[84] : level4[85];
	assign level5[43] = s[5] ? level4[86] : level4[87];
	assign level5[44] = s[5] ? level4[88] : level4[89];
	assign level5[45] = s[5] ? level4[90] : level4[91];
	assign level5[46] = s[5] ? level4[92] : level4[93];
	assign level5[47] = s[5] ? level4[94] : level4[95];
	assign level5[48] = s[5] ? level4[96] : level4[97];
	assign level5[49] = s[5] ? level4[98] : level4[99];
	assign level5[50] = s[5] ? level4[100] : level4[101];
	assign level5[51] = s[5] ? level4[102] : level4[103];
	assign level5[52] = s[5] ? level4[104] : level4[105];
	assign level5[53] = s[5] ? level4[106] : level4[107];
	assign level5[54] = s[5] ? level4[108] : level4[109];
	assign level5[55] = s[5] ? level4[110] : level4[111];
	assign level5[56] = s[5] ? level4[112] : level4[113];
	assign level5[57] = s[5] ? level4[114] : level4[115];
	assign level5[58] = s[5] ? level4[116] : level4[117];
	assign level5[59] = s[5] ? level4[118] : level4[119];
	assign level5[60] = s[5] ? level4[120] : level4[121];
	assign level5[61] = s[5] ? level4[122] : level4[123];
	assign level5[62] = s[5] ? level4[124] : level4[125];
	assign level5[63] = s[5] ? level4[126] : level4[127];

	assign level6[0] = s[6] ? level5[0] : level5[1];
	assign level6[1] = s[6] ? level5[2] : level5[3];
	assign level6[2] = s[6] ? level5[4] : level5[5];
	assign level6[3] = s[6] ? level5[6] : level5[7];
	assign level6[4] = s[6] ? level5[8] : level5[9];
	assign level6[5] = s[6] ? level5[10] : level5[11];
	assign level6[6] = s[6] ? level5[12] : level5[13];
	assign level6[7] = s[6] ? level5[14] : level5[15];
	assign level6[8] = s[6] ? level5[16] : level5[17];
	assign level6[9] = s[6] ? level5[18] : level5[19];
	assign level6[10] = s[6] ? level5[20] : level5[21];
	assign level6[11] = s[6] ? level5[22] : level5[23];
	assign level6[12] = s[6] ? level5[24] : level5[25];
	assign level6[13] = s[6] ? level5[26] : level5[27];
	assign level6[14] = s[6] ? level5[28] : level5[29];
	assign level6[15] = s[6] ? level5[30] : level5[31];
	assign level6[16] = s[6] ? level5[32] : level5[33];
	assign level6[17] = s[6] ? level5[34] : level5[35];
	assign level6[18] = s[6] ? level5[36] : level5[37];
	assign level6[19] = s[6] ? level5[38] : level5[39];
	assign level6[20] = s[6] ? level5[40] : level5[41];
	assign level6[21] = s[6] ? level5[42] : level5[43];
	assign level6[22] = s[6] ? level5[44] : level5[45];
	assign level6[23] = s[6] ? level5[46] : level5[47];
	assign level6[24] = s[6] ? level5[48] : level5[49];
	assign level6[25] = s[6] ? level5[50] : level5[51];
	assign level6[26] = s[6] ? level5[52] : level5[53];
	assign level6[27] = s[6] ? level5[54] : level5[55];
	assign level6[28] = s[6] ? level5[56] : level5[57];
	assign level6[29] = s[6] ? level5[58] : level5[59];
	assign level6[30] = s[6] ? level5[60] : level5[61];
	assign level6[31] = s[6] ? level5[62] : level5[63];

	assign level7[0] = s[7] ? level6[0] : level6[1];
	assign level7[1] = s[7] ? level6[2] : level6[3];
	assign level7[2] = s[7] ? level6[4] : level6[5];
	assign level7[3] = s[7] ? level6[6] : level6[7];
	assign level7[4] = s[7] ? level6[8] : level6[9];
	assign level7[5] = s[7] ? level6[10] : level6[11];
	assign level7[6] = s[7] ? level6[12] : level6[13];
	assign level7[7] = s[7] ? level6[14] : level6[15];
	assign level7[8] = s[7] ? level6[16] : level6[17];
	assign level7[9] = s[7] ? level6[18] : level6[19];
	assign level7[10] = s[7] ? level6[20] : level6[21];
	assign level7[11] = s[7] ? level6[22] : level6[23];
	assign level7[12] = s[7] ? level6[24] : level6[25];
	assign level7[13] = s[7] ? level6[26] : level6[27];
	assign level7[14] = s[7] ? level6[28] : level6[29];
	assign level7[15] = s[7] ? level6[30] : level6[31];

	assign level8[0] = s[8] ? level7[0] : level7[1];
	assign level8[1] = s[8] ? level7[2] : level7[3];
	assign level8[2] = s[8] ? level7[4] : level7[5];
	assign level8[3] = s[8] ? level7[6] : level7[7];
	assign level8[4] = s[8] ? level7[8] : level7[9];
	assign level8[5] = s[8] ? level7[10] : level7[11];
	assign level8[6] = s[8] ? level7[12] : level7[13];
	assign level8[7] = s[8] ? level7[14] : level7[15];

	assign level9[0] = s[9] ? level8[0] : level8[1];
	assign level9[1] = s[9] ? level8[2] : level8[3];
	assign level9[2] = s[9] ? level8[4] : level8[5];
	assign level9[3] = s[9] ? level8[6] : level8[7];

	assign level10[0] = s[10] ? level9[0] : level9[1];
	assign level10[1] = s[10] ? level9[2] : level9[3];

	assign level11[0] = s[11] ? level10[0] : level10[1];

	assign out = level11[0];
endmodule


module en_counter0 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


module en_counter1 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


module en_counter2 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


module en_counter3 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


module en_counter4 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


module en_counter5 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


module en_counter6 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


module en_counter7 (
	input  clock, reset,
	input  logic en,
	output logic [11:0] out
);
	always_ff @(posedge clock) begin
		if      (reset == 1)   out <= 'b0;
		else if (en == 1)      out <= out + 1;
		else                   out <= out - 1;
	end
endmodule


// Top level module
module filter (
	input  clock, reset,
	input  logic [11:0]  in,
	output logic [11:0]  outs [7:0]
);
	logic [11:0] pcc_in [148:0];
	logic       pos_SNs         [148:0];
	logic       neg_SNs         [148:0];
	logic [11:0] s;
	logic [11:0] r;
	logic       tree_outs [7:0];
	control crtl(.clock(clock), .reset(reset), .in(in), .out(pcc_in));
	counter cnt(.clock(clock), .reset(reset), .rev_state(r), .state(s));
	comparator_array_pos pccs_pos(.in(pcc_in), .r(r[11:0]), .xs(pos_SNs));
	comparator_array_neg pccs_neg(.in(pcc_in), .r(r[11:0]), .xs(neg_SNs));
	hw_tree0 tree0(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[0]));
	en_counter0 est0(.clock(clock), .reset(reset), .en(tree_outs[0]), .out(outs[0]));
	hw_tree1 tree1(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[1]));
	en_counter1 est1(.clock(clock), .reset(reset), .en(tree_outs[1]), .out(outs[1]));
	hw_tree2 tree2(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[2]));
	en_counter2 est2(.clock(clock), .reset(reset), .en(tree_outs[2]), .out(outs[2]));
	hw_tree3 tree3(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[3]));
	en_counter3 est3(.clock(clock), .reset(reset), .en(tree_outs[3]), .out(outs[3]));
	hw_tree4 tree4(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[4]));
	en_counter4 est4(.clock(clock), .reset(reset), .en(tree_outs[4]), .out(outs[4]));
	hw_tree5 tree5(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[5]));
	en_counter5 est5(.clock(clock), .reset(reset), .en(tree_outs[5]), .out(outs[5]));
	hw_tree6 tree6(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[6]));
	en_counter6 est6(.clock(clock), .reset(reset), .en(tree_outs[6]), .out(outs[6]));
	hw_tree7 tree7(.pos_SNs(pos_SNs), .neg_SNs(neg_SNs), .s(s), .out(tree_outs[7]));
	en_counter7 est7(.clock(clock), .reset(reset), .en(tree_outs[7]), .out(outs[7]));
endmodule