localparam [`len_idx-1:0] mapping[`pow2n-1:0] = {`len_idx'd0, `len_idx'd0, `len_idx'd0, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd2, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4,\
`len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd4, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6,\
`len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6,\
`len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6,\
`len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6,\
`len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd6, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8, `len_idx'd8,\
`len_idx'd8, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9,\
`len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd9, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10,\
`len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd10, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12,\
`len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12,\
`len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12,\
`len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12,\
`len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd12, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14,\
`len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd14, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd16, `len_idx'd18, `len_idx'd18, `len_idx'd18};