`define n 12
`define pow2n 4096
`define order 18
`define length 19
`define len_idx 5 // ceil(log2(19))=5
